`timescale 1 ns/100 ps
// Version: 


module MSS_075(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MGPIO0B_IN,
       MGPIO10B_IN,
       MGPIO1B_IN,
       MGPIO25A_IN,
       MGPIO26A_IN,
       MGPIO27A_IN,
       MGPIO28A_IN,
       MGPIO29A_IN,
       MGPIO2B_IN,
       MGPIO30A_IN,
       MGPIO31A_IN,
       MGPIO3B_IN,
       MGPIO4B_IN,
       MGPIO5B_IN,
       MGPIO6B_IN,
       MGPIO7B_IN,
       MGPIO8B_IN,
       MGPIO9B_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_CTS_MGPIO13B_IN,
       MMUART1_DCD_MGPIO16B_IN,
       MMUART1_DSR_MGPIO14B_IN,
       MMUART1_DTR_MGPIO12B_IN,
       MMUART1_RI_MGPIO15B_IN,
       MMUART1_RTS_MGPIO11B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI0_SS4_MGPIO19A_IN,
       SPI0_SS5_MGPIO20A_IN,
       SPI0_SS6_MGPIO21A_IN,
       SPI0_SS7_MGPIO22A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       USBD_DATA0_IN,
       USBD_DATA1_IN,
       USBD_DATA2_IN,
       USBD_DATA3_IN,
       USBD_DATA4_IN,
       USBD_DATA5_IN,
       USBD_DATA6_IN,
       USBD_DATA7_MGPIO23B_IN,
       USBD_DIR_IN,
       USBD_NXT_IN,
       USBD_STP_IN,
       USBD_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MGPIO0B_OUT,
       MGPIO10B_OUT,
       MGPIO1B_OUT,
       MGPIO25A_OUT,
       MGPIO26A_OUT,
       MGPIO27A_OUT,
       MGPIO28A_OUT,
       MGPIO29A_OUT,
       MGPIO2B_OUT,
       MGPIO30A_OUT,
       MGPIO31A_OUT,
       MGPIO3B_OUT,
       MGPIO4B_OUT,
       MGPIO5B_OUT,
       MGPIO6B_OUT,
       MGPIO7B_OUT,
       MGPIO8B_OUT,
       MGPIO9B_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_CTS_MGPIO13B_OUT,
       MMUART1_DCD_MGPIO16B_OUT,
       MMUART1_DSR_MGPIO14B_OUT,
       MMUART1_DTR_MGPIO12B_OUT,
       MMUART1_RI_MGPIO15B_OUT,
       MMUART1_RTS_MGPIO11B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI0_SS4_MGPIO19A_OUT,
       SPI0_SS5_MGPIO20A_OUT,
       SPI0_SS6_MGPIO21A_OUT,
       SPI0_SS7_MGPIO22A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       USBD_DATA0_OUT,
       USBD_DATA1_OUT,
       USBD_DATA2_OUT,
       USBD_DATA3_OUT,
       USBD_DATA4_OUT,
       USBD_DATA5_OUT,
       USBD_DATA6_OUT,
       USBD_DATA7_MGPIO23B_OUT,
       USBD_DIR_OUT,
       USBD_NXT_OUT,
       USBD_STP_OUT,
       USBD_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MGPIO0B_OE,
       MGPIO10B_OE,
       MGPIO1B_OE,
       MGPIO25A_OE,
       MGPIO26A_OE,
       MGPIO27A_OE,
       MGPIO28A_OE,
       MGPIO29A_OE,
       MGPIO2B_OE,
       MGPIO30A_OE,
       MGPIO31A_OE,
       MGPIO3B_OE,
       MGPIO4B_OE,
       MGPIO5B_OE,
       MGPIO6B_OE,
       MGPIO7B_OE,
       MGPIO8B_OE,
       MGPIO9B_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_CTS_MGPIO13B_OE,
       MMUART1_DCD_MGPIO16B_OE,
       MMUART1_DSR_MGPIO14B_OE,
       MMUART1_DTR_MGPIO12B_OE,
       MMUART1_RI_MGPIO15B_OE,
       MMUART1_RTS_MGPIO11B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI0_SS4_MGPIO19A_OE,
       SPI0_SS5_MGPIO20A_OE,
       SPI0_SS6_MGPIO21A_OE,
       SPI0_SS7_MGPIO22A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE,
       USBD_DATA0_OE,
       USBD_DATA1_OE,
       USBD_DATA2_OE,
       USBD_DATA3_OE,
       USBD_DATA4_OE,
       USBD_DATA5_OE,
       USBD_DATA6_OE,
       USBD_DATA7_MGPIO23B_OE,
       USBD_DIR_OE,
       USBD_NXT_OE,
       USBD_STP_OE,
       USBD_XCLK_OE
    ) ;
/* synthesis syn_black_box

syn_tsu0 = " CAN_RXBUS_F2H_SCP->CLK_BASE = 1.251"
syn_tsu1 = " F2HCALIB->CLK_BASE = 0.168"
syn_tsu2 = " F_FM0_ADDR[0]->CLK_BASE = 1.222"
syn_tsu3 = " F_FM0_ADDR[10]->CLK_BASE = 1.498"
syn_tsu4 = " F_FM0_ADDR[11]->CLK_BASE = 1.465"
syn_tsu5 = " F_FM0_ADDR[12]->CLK_BASE = 1.329"
syn_tsu6 = " F_FM0_ADDR[13]->CLK_BASE = 1.469"
syn_tsu7 = " F_FM0_ADDR[14]->CLK_BASE = 1.234"
syn_tsu8 = " F_FM0_ADDR[15]->CLK_BASE = 1.203"
syn_tsu9 = " F_FM0_ADDR[16]->CLK_BASE = 1.182"
syn_tsu10 = " F_FM0_ADDR[17]->CLK_BASE = 1.464"
syn_tsu11 = " F_FM0_ADDR[18]->CLK_BASE = 1.517"
syn_tsu12 = " F_FM0_ADDR[19]->CLK_BASE = 1.133"
syn_tsu13 = " F_FM0_ADDR[1]->CLK_BASE = 1.143"
syn_tsu14 = " F_FM0_ADDR[20]->CLK_BASE = 1.466"
syn_tsu15 = " F_FM0_ADDR[21]->CLK_BASE = 1.435"
syn_tsu16 = " F_FM0_ADDR[22]->CLK_BASE = 1.201"
syn_tsu17 = " F_FM0_ADDR[23]->CLK_BASE = 1.431"
syn_tsu18 = " F_FM0_ADDR[24]->CLK_BASE = 1.397"
syn_tsu19 = " F_FM0_ADDR[25]->CLK_BASE = 1.438"
syn_tsu20 = " F_FM0_ADDR[26]->CLK_BASE = 1.392"
syn_tsu21 = " F_FM0_ADDR[27]->CLK_BASE = 1.418"
syn_tsu22 = " F_FM0_ADDR[28]->CLK_BASE = 1.185"
syn_tsu23 = " F_FM0_ADDR[29]->CLK_BASE = 1.458"
syn_tsu24 = " F_FM0_ADDR[2]->CLK_BASE = 1.15"
syn_tsu25 = " F_FM0_ADDR[30]->CLK_BASE = 1.212"
syn_tsu26 = " F_FM0_ADDR[31]->CLK_BASE = 1.293"
syn_tsu27 = " F_FM0_ADDR[3]->CLK_BASE = 1.363"
syn_tsu28 = " F_FM0_ADDR[4]->CLK_BASE = 1.52"
syn_tsu29 = " F_FM0_ADDR[5]->CLK_BASE = 1.448"
syn_tsu30 = " F_FM0_ADDR[6]->CLK_BASE = 1.102"
syn_tsu31 = " F_FM0_ADDR[7]->CLK_BASE = 1.216"
syn_tsu32 = " F_FM0_ADDR[8]->CLK_BASE = 1.472"
syn_tsu33 = " F_FM0_ADDR[9]->CLK_BASE = 1.2"
syn_tsu34 = " F_FM0_ENABLE->CLK_BASE = 1.125"
syn_tsu35 = " F_FM0_SEL->CLK_BASE = 1.209"
syn_tsu36 = " F_FM0_WDATA[0]->CLK_BASE = 1.192"
syn_tsu37 = " F_FM0_WDATA[10]->CLK_BASE = 1.199"
syn_tsu38 = " F_FM0_WDATA[11]->CLK_BASE = 0.914"
syn_tsu39 = " F_FM0_WDATA[12]->CLK_BASE = 1.259"
syn_tsu40 = " F_FM0_WDATA[13]->CLK_BASE = 0.343"
syn_tsu41 = " F_FM0_WDATA[14]->CLK_BASE = 1.23"
syn_tsu42 = " F_FM0_WDATA[15]->CLK_BASE = 1.314"
syn_tsu43 = " F_FM0_WDATA[16]->CLK_BASE = 1.186"
syn_tsu44 = " F_FM0_WDATA[17]->CLK_BASE = 1.185"
syn_tsu45 = " F_FM0_WDATA[18]->CLK_BASE = 1.232"
syn_tsu46 = " F_FM0_WDATA[19]->CLK_BASE = 1.213"
syn_tsu47 = " F_FM0_WDATA[1]->CLK_BASE = 1.327"
syn_tsu48 = " F_FM0_WDATA[20]->CLK_BASE = 1.248"
syn_tsu49 = " F_FM0_WDATA[21]->CLK_BASE = 1.135"
syn_tsu50 = " F_FM0_WDATA[22]->CLK_BASE = 1.201"
syn_tsu51 = " F_FM0_WDATA[23]->CLK_BASE = 1.217"
syn_tsu52 = " F_FM0_WDATA[24]->CLK_BASE = 1.193"
syn_tsu53 = " F_FM0_WDATA[25]->CLK_BASE = 1.251"
syn_tsu54 = " F_FM0_WDATA[26]->CLK_BASE = 1.211"
syn_tsu55 = " F_FM0_WDATA[27]->CLK_BASE = 1.155"
syn_tsu56 = " F_FM0_WDATA[28]->CLK_BASE = 1.185"
syn_tsu57 = " F_FM0_WDATA[29]->CLK_BASE = 1.156"
syn_tsu58 = " F_FM0_WDATA[2]->CLK_BASE = 0.947"
syn_tsu59 = " F_FM0_WDATA[30]->CLK_BASE = 1.24"
syn_tsu60 = " F_FM0_WDATA[31]->CLK_BASE = 1.194"
syn_tsu61 = " F_FM0_WDATA[3]->CLK_BASE = 1.253"
syn_tsu62 = " F_FM0_WDATA[4]->CLK_BASE = 1.252"
syn_tsu63 = " F_FM0_WDATA[5]->CLK_BASE = 1.272"
syn_tsu64 = " F_FM0_WDATA[6]->CLK_BASE = 1.205"
syn_tsu65 = " F_FM0_WDATA[7]->CLK_BASE = 1.285"
syn_tsu66 = " F_FM0_WDATA[8]->CLK_BASE = 1.182"
syn_tsu67 = " F_FM0_WDATA[9]->CLK_BASE = 1.181"
syn_tsu68 = " F_FM0_WRITE->CLK_BASE = 1.137"
syn_tsu69 = " F_HM0_RDATA[0]->CLK_BASE = 0.964"
syn_tsu70 = " F_HM0_RDATA[10]->CLK_BASE = 0.974"
syn_tsu71 = " F_HM0_RDATA[11]->CLK_BASE = 0.98"
syn_tsu72 = " F_HM0_RDATA[12]->CLK_BASE = 0.991"
syn_tsu73 = " F_HM0_RDATA[13]->CLK_BASE = 1.107"
syn_tsu74 = " F_HM0_RDATA[14]->CLK_BASE = 1.067"
syn_tsu75 = " F_HM0_RDATA[15]->CLK_BASE = 1.09"
syn_tsu76 = " F_HM0_RDATA[16]->CLK_BASE = 1.059"
syn_tsu77 = " F_HM0_RDATA[17]->CLK_BASE = 1.185"
syn_tsu78 = " F_HM0_RDATA[18]->CLK_BASE = 1.282"
syn_tsu79 = " F_HM0_RDATA[19]->CLK_BASE = 1.105"
syn_tsu80 = " F_HM0_RDATA[1]->CLK_BASE = 1.015"
syn_tsu81 = " F_HM0_RDATA[20]->CLK_BASE = 1.096"
syn_tsu82 = " F_HM0_RDATA[21]->CLK_BASE = 1.136"
syn_tsu83 = " F_HM0_RDATA[22]->CLK_BASE = 1.355"
syn_tsu84 = " F_HM0_RDATA[23]->CLK_BASE = 1.104"
syn_tsu85 = " F_HM0_RDATA[24]->CLK_BASE = 1.04"
syn_tsu86 = " F_HM0_RDATA[25]->CLK_BASE = 1.098"
syn_tsu87 = " F_HM0_RDATA[26]->CLK_BASE = 1.151"
syn_tsu88 = " F_HM0_RDATA[27]->CLK_BASE = 1.1"
syn_tsu89 = " F_HM0_RDATA[28]->CLK_BASE = 1.115"
syn_tsu90 = " F_HM0_RDATA[29]->CLK_BASE = 1.158"
syn_tsu91 = " F_HM0_RDATA[2]->CLK_BASE = 1.297"
syn_tsu92 = " F_HM0_RDATA[30]->CLK_BASE = 1.161"
syn_tsu93 = " F_HM0_RDATA[31]->CLK_BASE = 1.051"
syn_tsu94 = " F_HM0_RDATA[3]->CLK_BASE = 0.955"
syn_tsu95 = " F_HM0_RDATA[4]->CLK_BASE = 0.99"
syn_tsu96 = " F_HM0_RDATA[5]->CLK_BASE = 0.976"
syn_tsu97 = " F_HM0_RDATA[6]->CLK_BASE = 0.947"
syn_tsu98 = " F_HM0_RDATA[7]->CLK_BASE = 1"
syn_tsu99 = " F_HM0_RDATA[8]->CLK_BASE = 0.995"
syn_tsu100 = " F_HM0_RDATA[9]->CLK_BASE = 1.034"
syn_tsu101 = " F_HM0_READY->CLK_BASE = 1.057"
syn_tsu102 = " F_HM0_RESP->CLK_BASE = 1.114"
syn_tsu103 = " I2C0_SDA_F2H_SCP->I2C0_SCL_F2H_SCP = 0.013"
syn_tsu104 = " I2C1_SDA_F2H_SCP->I2C1_SCL_F2H_SCP = 0.255"
syn_tsu105 = " MGPIO0A_F2H_GPIN->CLK_BASE = 0.251"
syn_tsu106 = " MGPIO10A_F2H_GPIN->CLK_BASE = 0.485"
syn_tsu107 = " MGPIO11A_F2H_GPIN->CLK_BASE = 0.469"
syn_tsu108 = " MGPIO11B_F2H_GPIN->CLK_BASE = 0.827"
syn_tsu109 = " MGPIO12A_F2H_GPIN->CLK_BASE = 0.485"
syn_tsu110 = " MGPIO13A_F2H_GPIN->CLK_BASE = 0.337"
syn_tsu111 = " MGPIO14A_F2H_GPIN->CLK_BASE = 0.355"
syn_tsu112 = " MGPIO15A_F2H_GPIN->CLK_BASE = 0.216"
syn_tsu113 = " MGPIO16A_F2H_GPIN->CLK_BASE = 0.35"
syn_tsu114 = " MGPIO17B_F2H_GPIN->CLK_BASE = 0.272"
syn_tsu115 = " MGPIO18B_F2H_GPIN->CLK_BASE = 0.273"
syn_tsu116 = " MGPIO19B_F2H_GPIN->CLK_BASE = 0.553"
syn_tsu117 = " MGPIO1A_F2H_GPIN->CLK_BASE = 0.388"
syn_tsu118 = " MGPIO20B_F2H_GPIN->CLK_BASE = 0.508"
syn_tsu119 = " MGPIO21B_F2H_GPIN->CLK_BASE = 0.261"
syn_tsu120 = " MGPIO22B_F2H_GPIN->CLK_BASE = 0.509"
syn_tsu121 = " MGPIO24B_F2H_GPIN->CLK_BASE = 0.515"
syn_tsu122 = " MGPIO25B_F2H_GPIN->CLK_BASE = 0.464"
syn_tsu123 = " MGPIO26B_F2H_GPIN->CLK_BASE = 0.516"
syn_tsu124 = " MGPIO27B_F2H_GPIN->CLK_BASE = 0.547"
syn_tsu125 = " MGPIO28B_F2H_GPIN->CLK_BASE = 0.642"
syn_tsu126 = " MGPIO29B_F2H_GPIN->CLK_BASE = 0.543"
syn_tsu127 = " MGPIO2A_F2H_GPIN->CLK_BASE = 0.188"
syn_tsu128 = " MGPIO30B_F2H_GPIN->CLK_BASE = 0.393"
syn_tsu129 = " MGPIO31B_F2H_GPIN->CLK_BASE = 0.496"
syn_tsu130 = " MGPIO3A_F2H_GPIN->CLK_BASE = 0.138"
syn_tsu131 = " MGPIO4A_F2H_GPIN->CLK_BASE = 0.257"
syn_tsu132 = " MGPIO5A_F2H_GPIN->CLK_BASE = 0.176"
syn_tsu133 = " MGPIO6A_F2H_GPIN->CLK_BASE = 0.246"
syn_tsu134 = " MGPIO7A_F2H_GPIN->CLK_BASE = 0.23"
syn_tsu135 = " MGPIO8A_F2H_GPIN->CLK_BASE = 0.353"
syn_tsu136 = " MGPIO9A_F2H_GPIN->CLK_BASE = 0.262"
syn_tsu137 = " MMUART0_CTS_F2H_SCP->CLK_BASE = 0.702"
syn_tsu138 = " MMUART0_DCD_F2H_SCP->CLK_BASE = 0.66"
syn_tsu139 = " MMUART0_DSR_F2H_SCP->CLK_BASE = 0.627"
syn_tsu140 = " MMUART0_RI_F2H_SCP->CLK_BASE = 0.557"
syn_tsu141 = " MMUART0_SCK_F2H_SCP->CLK_BASE = 0.284"
syn_tsu142 = " MMUART0_TXD_F2H_SCP->CLK_BASE = 0.656"
syn_tsu143 = " MMUART1_CTS_F2H_SCP->CLK_BASE = 1.03"
syn_tsu144 = " MMUART1_DCD_F2H_SCP->CLK_BASE = 0.636"
syn_tsu145 = " MMUART1_DSR_F2H_SCP->CLK_BASE = 0.825"
syn_tsu146 = " MMUART1_RI_F2H_SCP->CLK_BASE = 0.566"
syn_tsu147 = " MMUART1_RXD_F2H_SCP->CLK_BASE = 0.842"
syn_tsu148 = " MMUART1_SCK_F2H_SCP->CLK_BASE = 0.859"
syn_tsu149 = " MMUART1_TXD_F2H_SCP->CLK_BASE = 0.806"
syn_tsu150 = " SMBALERT_NI0->I2C0_SCL_F2H_SCP = 0"
syn_tsu151 = " SMBALERT_NI1->I2C1_SCL_F2H_SCP = 0"
syn_tsu152 = " SMBSUS_NI0->I2C0_SCL_F2H_SCP = 0"
syn_tsu153 = " SMBSUS_NI1->I2C1_SCL_F2H_SCP = 0"
syn_tsu154 = " SPI1_SDI_F2H_SCP->SPI1_CLK_IN = 0.617"
syn_tco0 = " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_A = 3.279"
syn_tco1 = " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_B = 2.868"
syn_tco2 = " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_A = 2.961"
syn_tco3 = " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_B = 2.973"
syn_tco4 = " CLK_BASE->CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT = 4.722"
syn_tco5 = " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_A = 2.884"
syn_tco6 = " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_B = 2.882"
syn_tco7 = " CLK_BASE->CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT = 4.447"
syn_tco8 = " CLK_BASE->F_FM0_RDATA[0] = 3.961"
syn_tco9 = " CLK_BASE->F_FM0_RDATA[10] = 3.977"
syn_tco10 = " CLK_BASE->F_FM0_RDATA[11] = 3.941"
syn_tco11 = " CLK_BASE->F_FM0_RDATA[12] = 3.884"
syn_tco12 = " CLK_BASE->F_FM0_RDATA[13] = 3.899"
syn_tco13 = " CLK_BASE->F_FM0_RDATA[14] = 3.926"
syn_tco14 = " CLK_BASE->F_FM0_RDATA[15] = 3.870"
syn_tco15 = " CLK_BASE->F_FM0_RDATA[16] = 3.686"
syn_tco16 = " CLK_BASE->F_FM0_RDATA[17] = 3.688"
syn_tco17 = " CLK_BASE->F_FM0_RDATA[18] = 3.719"
syn_tco18 = " CLK_BASE->F_FM0_RDATA[19] = 3.577"
syn_tco19 = " CLK_BASE->F_FM0_RDATA[1] = 3.932"
syn_tco20 = " CLK_BASE->F_FM0_RDATA[20] = 3.614"
syn_tco21 = " CLK_BASE->F_FM0_RDATA[21] = 3.600"
syn_tco22 = " CLK_BASE->F_FM0_RDATA[22] = 3.737"
syn_tco23 = " CLK_BASE->F_FM0_RDATA[23] = 3.681"
syn_tco24 = " CLK_BASE->F_FM0_RDATA[24] = 3.605"
syn_tco25 = " CLK_BASE->F_FM0_RDATA[25] = 3.590"
syn_tco26 = " CLK_BASE->F_FM0_RDATA[26] = 3.680"
syn_tco27 = " CLK_BASE->F_FM0_RDATA[27] = 3.703"
syn_tco28 = " CLK_BASE->F_FM0_RDATA[28] = 3.707"
syn_tco29 = " CLK_BASE->F_FM0_RDATA[29] = 3.696"
syn_tco30 = " CLK_BASE->F_FM0_RDATA[2] = 3.916"
syn_tco31 = " CLK_BASE->F_FM0_RDATA[30] = 3.669"
syn_tco32 = " CLK_BASE->F_FM0_RDATA[31] = 3.585"
syn_tco33 = " CLK_BASE->F_FM0_RDATA[3] = 3.908"
syn_tco34 = " CLK_BASE->F_FM0_RDATA[4] = 3.986"
syn_tco35 = " CLK_BASE->F_FM0_RDATA[5] = 3.941"
syn_tco36 = " CLK_BASE->F_FM0_RDATA[6] = 3.897"
syn_tco37 = " CLK_BASE->F_FM0_RDATA[7] = 3.924"
syn_tco38 = " CLK_BASE->F_FM0_RDATA[8] = 3.912"
syn_tco39 = " CLK_BASE->F_FM0_RDATA[9] = 3.938"
syn_tco40 = " CLK_BASE->F_FM0_READYOUT = 3.443"
syn_tco41 = " CLK_BASE->F_FM0_RESP = 3.356"
syn_tco42 = " CLK_BASE->F_HM0_ADDR[0] = 3.056"
syn_tco43 = " CLK_BASE->F_HM0_ADDR[10] = 3.153"
syn_tco44 = " CLK_BASE->F_HM0_ADDR[11] = 3.035"
syn_tco45 = " CLK_BASE->F_HM0_ADDR[12] = 3.046"
syn_tco46 = " CLK_BASE->F_HM0_ADDR[13] = 3.017"
syn_tco47 = " CLK_BASE->F_HM0_ADDR[14] = 3.012"
syn_tco48 = " CLK_BASE->F_HM0_ADDR[15] = 3.056"
syn_tco49 = " CLK_BASE->F_HM0_ADDR[16] = 3.101"
syn_tco50 = " CLK_BASE->F_HM0_ADDR[17] = 3.126"
syn_tco51 = " CLK_BASE->F_HM0_ADDR[18] = 3.114"
syn_tco52 = " CLK_BASE->F_HM0_ADDR[19] = 3.116"
syn_tco53 = " CLK_BASE->F_HM0_ADDR[1] = 3.038"
syn_tco54 = " CLK_BASE->F_HM0_ADDR[20] = 3.146"
syn_tco55 = " CLK_BASE->F_HM0_ADDR[21] = 3.034"
syn_tco56 = " CLK_BASE->F_HM0_ADDR[22] = 3.006"
syn_tco57 = " CLK_BASE->F_HM0_ADDR[23] = 3.052"
syn_tco58 = " CLK_BASE->F_HM0_ADDR[24] = 3.023"
syn_tco59 = " CLK_BASE->F_HM0_ADDR[25] = 3.051"
syn_tco60 = " CLK_BASE->F_HM0_ADDR[26] = 3.053"
syn_tco61 = " CLK_BASE->F_HM0_ADDR[27] = 3.030"
syn_tco62 = " CLK_BASE->F_HM0_ADDR[28] = 3.022"
syn_tco63 = " CLK_BASE->F_HM0_ADDR[29] = 3.020"
syn_tco64 = " CLK_BASE->F_HM0_ADDR[2] = 3.014"
syn_tco65 = " CLK_BASE->F_HM0_ADDR[30] = 3.018"
syn_tco66 = " CLK_BASE->F_HM0_ADDR[31] = 3.031"
syn_tco67 = " CLK_BASE->F_HM0_ADDR[3] = 3.035"
syn_tco68 = " CLK_BASE->F_HM0_ADDR[4] = 3.187"
syn_tco69 = " CLK_BASE->F_HM0_ADDR[5] = 3.021"
syn_tco70 = " CLK_BASE->F_HM0_ADDR[6] = 3.131"
syn_tco71 = " CLK_BASE->F_HM0_ADDR[7] = 3.033"
syn_tco72 = " CLK_BASE->F_HM0_ADDR[8] = 3.128"
syn_tco73 = " CLK_BASE->F_HM0_ADDR[9] = 3.042"
syn_tco74 = " CLK_BASE->F_HM0_ENABLE = 3.250"
syn_tco75 = " CLK_BASE->F_HM0_SEL = 3.083"
syn_tco76 = " CLK_BASE->F_HM0_WDATA[0] = 3.205"
syn_tco77 = " CLK_BASE->F_HM0_WDATA[10] = 3.059"
syn_tco78 = " CLK_BASE->F_HM0_WDATA[11] = 3.078"
syn_tco79 = " CLK_BASE->F_HM0_WDATA[12] = 3.067"
syn_tco80 = " CLK_BASE->F_HM0_WDATA[13] = 3.067"
syn_tco81 = " CLK_BASE->F_HM0_WDATA[14] = 3.079"
syn_tco82 = " CLK_BASE->F_HM0_WDATA[15] = 3.081"
syn_tco83 = " CLK_BASE->F_HM0_WDATA[16] = 3.063"
syn_tco84 = " CLK_BASE->F_HM0_WDATA[17] = 3.042"
syn_tco85 = " CLK_BASE->F_HM0_WDATA[18] = 3.069"
syn_tco86 = " CLK_BASE->F_HM0_WDATA[19] = 3.057"
syn_tco87 = " CLK_BASE->F_HM0_WDATA[1] = 3.180"
syn_tco88 = " CLK_BASE->F_HM0_WDATA[20] = 3.066"
syn_tco89 = " CLK_BASE->F_HM0_WDATA[21] = 3.055"
syn_tco90 = " CLK_BASE->F_HM0_WDATA[22] = 3.041"
syn_tco91 = " CLK_BASE->F_HM0_WDATA[23] = 3.057"
syn_tco92 = " CLK_BASE->F_HM0_WDATA[24] = 3.051"
syn_tco93 = " CLK_BASE->F_HM0_WDATA[25] = 3.029"
syn_tco94 = " CLK_BASE->F_HM0_WDATA[26] = 3.034"
syn_tco95 = " CLK_BASE->F_HM0_WDATA[27] = 3.024"
syn_tco96 = " CLK_BASE->F_HM0_WDATA[28] = 3.073"
syn_tco97 = " CLK_BASE->F_HM0_WDATA[29] = 3.065"
syn_tco98 = " CLK_BASE->F_HM0_WDATA[2] = 3.224"
syn_tco99 = " CLK_BASE->F_HM0_WDATA[30] = 3.030"
syn_tco100 = " CLK_BASE->F_HM0_WDATA[31] = 3.030"
syn_tco101 = " CLK_BASE->F_HM0_WDATA[3] = 3.171"
syn_tco102 = " CLK_BASE->F_HM0_WDATA[4] = 3.082"
syn_tco103 = " CLK_BASE->F_HM0_WDATA[5] = 3.085"
syn_tco104 = " CLK_BASE->F_HM0_WDATA[6] = 3.087"
syn_tco105 = " CLK_BASE->F_HM0_WDATA[7] = 3.078"
syn_tco106 = " CLK_BASE->F_HM0_WDATA[8] = 3.093"
syn_tco107 = " CLK_BASE->F_HM0_WDATA[9] = 3.083"
syn_tco108 = " CLK_BASE->F_HM0_WRITE = 3.119"
syn_tco109 = " CLK_BASE->H2FCALIB = 3.142"
syn_tco110 = " CLK_BASE->I2C0_SCL_MGPIO31B_H2F_B = 3.199"
syn_tco111 = " CLK_BASE->I2C0_SCL_USBC_DATA1_MGPIO31B_OE = 2.905"
syn_tco112 = " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_A = 3.052"
syn_tco113 = " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_B = 3.114"
syn_tco114 = " CLK_BASE->I2C0_SDA_USBC_DATA0_MGPIO30B_OE = 2.477"
syn_tco115 = " CLK_BASE->I2C1_SCL_MGPIO1A_H2F_B = 3.195"
syn_tco116 = " CLK_BASE->I2C1_SCL_USBA_DATA4_MGPIO1A_OE = 3.478"
syn_tco117 = " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_A = 2.807"
syn_tco118 = " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_B = 3.208"
syn_tco119 = " CLK_BASE->I2C1_SDA_USBA_DATA3_MGPIO0A_OE = 3.249"
syn_tco120 = " CLK_BASE->MGPIO0B_OE = 2.385"
syn_tco121 = " CLK_BASE->MGPIO0B_OUT = 2.393"
syn_tco122 = " CLK_BASE->MGPIO10B_OE = 2.180"
syn_tco123 = " CLK_BASE->MGPIO10B_OUT = 2.172"
syn_tco124 = " CLK_BASE->MGPIO1B_OE = 2.379"
syn_tco125 = " CLK_BASE->MGPIO1B_OUT = 2.487"
syn_tco126 = " CLK_BASE->MGPIO25A_OE = 4.208"
syn_tco127 = " CLK_BASE->MGPIO25A_OUT = 3.932"
syn_tco128 = " CLK_BASE->MGPIO26A_OE = 4.030"
syn_tco129 = " CLK_BASE->MGPIO26A_OUT = 4.008"
syn_tco130 = " CLK_BASE->MGPIO27A_OE = 3.746"
syn_tco131 = " CLK_BASE->MGPIO27A_OUT = 3.785"
syn_tco132 = " CLK_BASE->MGPIO28A_OE = 3.854"
syn_tco133 = " CLK_BASE->MGPIO28A_OUT = 4.121"
syn_tco134 = " CLK_BASE->MGPIO29A_OE = 2.439"
syn_tco135 = " CLK_BASE->MGPIO29A_OUT = 2.657"
syn_tco136 = " CLK_BASE->MGPIO2B_OE = 2.572"
syn_tco137 = " CLK_BASE->MGPIO2B_OUT = 2.430"
syn_tco138 = " CLK_BASE->MGPIO30A_OE = 2.652"
syn_tco139 = " CLK_BASE->MGPIO30A_OUT = 2.467"
syn_tco140 = " CLK_BASE->MGPIO31A_OE = 2.504"
syn_tco141 = " CLK_BASE->MGPIO31A_OUT = 2.581"
syn_tco142 = " CLK_BASE->MGPIO3B_OE = 2.384"
syn_tco143 = " CLK_BASE->MGPIO3B_OUT = 2.583"
syn_tco144 = " CLK_BASE->MGPIO4B_OE = 2.485"
syn_tco145 = " CLK_BASE->MGPIO4B_OUT = 2.270"
syn_tco146 = " CLK_BASE->MGPIO5B_OE = 2.601"
syn_tco147 = " CLK_BASE->MGPIO5B_OUT = 2.563"
syn_tco148 = " CLK_BASE->MGPIO6B_OE = 2.248"
syn_tco149 = " CLK_BASE->MGPIO6B_OUT = 2.364"
syn_tco150 = " CLK_BASE->MGPIO7B_OE = 2.273"
syn_tco151 = " CLK_BASE->MGPIO7B_OUT = 2.511"
syn_tco152 = " CLK_BASE->MGPIO8B_OE = 2.407"
syn_tco153 = " CLK_BASE->MGPIO8B_OUT = 2.398"
syn_tco154 = " CLK_BASE->MGPIO9B_OE = 2.228"
syn_tco155 = " CLK_BASE->MGPIO9B_OUT = 2.108"
syn_tco156 = " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_A = 3.124"
syn_tco157 = " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_B = 3.308"
syn_tco158 = " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_A = 3.025"
syn_tco159 = " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_B = 2.910"
syn_tco160 = " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_A = 3.289"
syn_tco161 = " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_B = 3.143"
syn_tco162 = " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_A = 2.850"
syn_tco163 = " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_B = 3.013"
syn_tco164 = " CLK_BASE->MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT = 2.489"
syn_tco165 = " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_A = 2.915"
syn_tco166 = " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_B = 2.882"
syn_tco167 = " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_A = 2.824"
syn_tco168 = " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_B = 2.958"
syn_tco169 = " CLK_BASE->MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT = 2.390"
syn_tco170 = " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_A = 3.026"
syn_tco171 = " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_B = 3.179"
syn_tco172 = " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_A = 3.146"
syn_tco173 = " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_B = 3.068"
syn_tco174 = " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OE = 2.799"
syn_tco175 = " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OUT = 2.265"
syn_tco176 = " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_A = 3.104"
syn_tco177 = " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_B = 3.227"
syn_tco178 = " CLK_BASE->MMUART0_TXD_USBC_DIR_MGPIO27B_OUT = 2.675"
syn_tco179 = " CLK_BASE->MMUART1_DTR_MGPIO12B_H2F_A = 3.201"
syn_tco180 = " CLK_BASE->MMUART1_DTR_MGPIO12B_OUT = 2.854"
syn_tco181 = " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_A = 3.148"
syn_tco182 = " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_B = 3.033"
syn_tco183 = " CLK_BASE->MMUART1_RTS_MGPIO11B_OUT = 3.209"
syn_tco184 = " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_A = 3.118"
syn_tco185 = " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_B = 3.235"
syn_tco186 = " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_A = 3.549"
syn_tco187 = " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_B = 3.424"
syn_tco188 = " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OE = 3.415"
syn_tco189 = " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT = 3.015"
syn_tco190 = " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_A = 3.024"
syn_tco191 = " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_B = 3.070"
syn_tco192 = " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OE = 3.510"
syn_tco193 = " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT = 3.004"
syn_tco194 = " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE = 4.835"
syn_tco195 = " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT = 4.518"
syn_tco196 = " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_A = 2.850"
syn_tco197 = " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_B = 3.216"
syn_tco198 = " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_A = 3.418"
syn_tco199 = " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_B = 2.942"
syn_tco200 = " CLK_BASE->SPI0_SDO_USBA_STP_MGPIO6A_OUT = 4.909"
syn_tco201 = " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_A = 3.312"
syn_tco202 = " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_B = 3.178"
syn_tco203 = " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_A = 3.277"
syn_tco204 = " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_B = 2.933"
syn_tco205 = " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_A = 3.370"
syn_tco206 = " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_B = 3.014"
syn_tco207 = " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_A = 3.333"
syn_tco208 = " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_B = 2.852"
syn_tco209 = " CLK_BASE->SPI0_SS4_MGPIO19A_H2F_A = 3.140"
syn_tco210 = " CLK_BASE->SPI0_SS5_MGPIO20A_H2F_A = 3.090"
syn_tco211 = " CLK_BASE->SPI0_SS6_MGPIO21A_H2F_A = 3.115"
syn_tco212 = " CLK_BASE->SPI0_SS7_MGPIO22A_H2F_A = 2.810"
syn_tco213 = " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_A = 3.365"
syn_tco214 = " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_B = 2.958"
syn_tco215 = " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_A = 3.179"
syn_tco216 = " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_B = 3.276"
syn_tco217 = " CLK_BASE->SPI1_SDO_MGPIO12A_OE = 5.662"
syn_tco218 = " CLK_BASE->SPI1_SDO_MGPIO12A_OUT = 5.344"
syn_tco219 = " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_A = 3.120"
syn_tco220 = " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_B = 3.102"
syn_tco221 = " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_A = 3.146"
syn_tco222 = " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_B = 3.343"
syn_tco223 = " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_A = 2.796"
syn_tco224 = " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_B = 2.794"
syn_tco225 = " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_A = 2.709"
syn_tco226 = " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_B = 3.367"
syn_tco227 = " CLK_BASE->SPI1_SS4_MGPIO17A_H2F_A = 2.916"
syn_tco228 = " CLK_BASE->SPI1_SS5_MGPIO18A_H2F_A = 2.933"
syn_tco229 = " CLK_BASE->SPI1_SS6_MGPIO23A_H2F_A = 3.008"
syn_tco230 = " CLK_BASE->SPI1_SS7_MGPIO24A_H2F_A = 2.971"
*/
/* synthesis black_box_pad_pin ="" */
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MGPIO0B_IN;
input  MGPIO10B_IN;
input  MGPIO1B_IN;
input  MGPIO25A_IN;
input  MGPIO26A_IN;
input  MGPIO27A_IN;
input  MGPIO28A_IN;
input  MGPIO29A_IN;
input  MGPIO2B_IN;
input  MGPIO30A_IN;
input  MGPIO31A_IN;
input  MGPIO3B_IN;
input  MGPIO4B_IN;
input  MGPIO5B_IN;
input  MGPIO6B_IN;
input  MGPIO7B_IN;
input  MGPIO8B_IN;
input  MGPIO9B_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_CTS_MGPIO13B_IN;
input  MMUART1_DCD_MGPIO16B_IN;
input  MMUART1_DSR_MGPIO14B_IN;
input  MMUART1_DTR_MGPIO12B_IN;
input  MMUART1_RI_MGPIO15B_IN;
input  MMUART1_RTS_MGPIO11B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI0_SS4_MGPIO19A_IN;
input  SPI0_SS5_MGPIO20A_IN;
input  SPI0_SS6_MGPIO21A_IN;
input  SPI0_SS7_MGPIO22A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
input  USBD_DATA0_IN;
input  USBD_DATA1_IN;
input  USBD_DATA2_IN;
input  USBD_DATA3_IN;
input  USBD_DATA4_IN;
input  USBD_DATA5_IN;
input  USBD_DATA6_IN;
input  USBD_DATA7_MGPIO23B_IN;
input  USBD_DIR_IN;
input  USBD_NXT_IN;
input  USBD_STP_IN;
input  USBD_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MGPIO0B_OUT;
output MGPIO10B_OUT;
output MGPIO1B_OUT;
output MGPIO25A_OUT;
output MGPIO26A_OUT;
output MGPIO27A_OUT;
output MGPIO28A_OUT;
output MGPIO29A_OUT;
output MGPIO2B_OUT;
output MGPIO30A_OUT;
output MGPIO31A_OUT;
output MGPIO3B_OUT;
output MGPIO4B_OUT;
output MGPIO5B_OUT;
output MGPIO6B_OUT;
output MGPIO7B_OUT;
output MGPIO8B_OUT;
output MGPIO9B_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_CTS_MGPIO13B_OUT;
output MMUART1_DCD_MGPIO16B_OUT;
output MMUART1_DSR_MGPIO14B_OUT;
output MMUART1_DTR_MGPIO12B_OUT;
output MMUART1_RI_MGPIO15B_OUT;
output MMUART1_RTS_MGPIO11B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI0_SS4_MGPIO19A_OUT;
output SPI0_SS5_MGPIO20A_OUT;
output SPI0_SS6_MGPIO21A_OUT;
output SPI0_SS7_MGPIO22A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output USBD_DATA0_OUT;
output USBD_DATA1_OUT;
output USBD_DATA2_OUT;
output USBD_DATA3_OUT;
output USBD_DATA4_OUT;
output USBD_DATA5_OUT;
output USBD_DATA6_OUT;
output USBD_DATA7_MGPIO23B_OUT;
output USBD_DIR_OUT;
output USBD_NXT_OUT;
output USBD_STP_OUT;
output USBD_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MGPIO0B_OE;
output MGPIO10B_OE;
output MGPIO1B_OE;
output MGPIO25A_OE;
output MGPIO26A_OE;
output MGPIO27A_OE;
output MGPIO28A_OE;
output MGPIO29A_OE;
output MGPIO2B_OE;
output MGPIO30A_OE;
output MGPIO31A_OE;
output MGPIO3B_OE;
output MGPIO4B_OE;
output MGPIO5B_OE;
output MGPIO6B_OE;
output MGPIO7B_OE;
output MGPIO8B_OE;
output MGPIO9B_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_CTS_MGPIO13B_OE;
output MMUART1_DCD_MGPIO16B_OE;
output MMUART1_DSR_MGPIO14B_OE;
output MMUART1_DTR_MGPIO12B_OE;
output MMUART1_RI_MGPIO15B_OE;
output MMUART1_RTS_MGPIO11B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI0_SS4_MGPIO19A_OE;
output SPI0_SS5_MGPIO20A_OE;
output SPI0_SS6_MGPIO21A_OE;
output SPI0_SS7_MGPIO22A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;
output USBD_DATA0_OE;
output USBD_DATA1_OE;
output USBD_DATA2_OE;
output USBD_DATA3_OE;
output USBD_DATA4_OE;
output USBD_DATA5_OE;
output USBD_DATA6_OE;
output USBD_DATA7_MGPIO23B_OE;
output USBD_DIR_OE;
output USBD_NXT_OE;
output USBD_STP_OE;
output USBD_XCLK_OE;
parameter INIT = 'h0;
parameter ACT_UBITS = 'h0;
parameter MEMORYFILE = "";
parameter RTC_MAIN_XTL_FREQ = 0.0;
parameter RTC_MAIN_XTL_MODE = "";
parameter DDR_CLK_FREQ = 0.0;

endmodule
