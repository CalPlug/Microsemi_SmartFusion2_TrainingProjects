`timescale 1 ns/100 ps
// Version: v11.7 11.7.0.119


module SERDESIF_075(
       APB_PRDATA,
       APB_PREADY,
       APB_PSLVERR,
       ATXCLKSTABLE,
       EPCS_READY,
       EPCS_RXCLK,
       EPCS_RXCLK_0,
       EPCS_RXCLK_1,
       EPCS_RXDATA,
       EPCS_RXIDLE,
       EPCS_RXRSTN,
       EPCS_RXVAL,
       EPCS_TXCLK,
       EPCS_TXCLK_0,
       EPCS_TXCLK_1,
       EPCS_TXRSTN,
       FATC_RESET_N,
       H2FCALIB0,
       H2FCALIB1,
       M2_ARADDR,
       M2_ARBURST,
       M2_ARID,
       M2_ARLEN,
       M2_ARSIZE,
       M2_ARVALID,
       M2_AWADDR_HADDR,
       M2_AWBURST_HTRANS,
       M2_AWID,
       M2_AWLEN_HBURST,
       M2_AWSIZE_HSIZE,
       M2_AWVALID_HWRITE,
       M2_BREADY,
       M2_RREADY,
       M2_WDATA_HWDATA,
       M2_WID,
       M2_WLAST,
       M2_WSTRB,
       M2_WVALID,
       M_ARADDR,
       M_ARBURST,
       M_ARID,
       M_ARLEN,
       M_ARSIZE,
       M_ARVALID,
       M_AWADDR_HADDR,
       M_AWBURST_HTRANS,
       M_AWID,
       M_AWLEN_HBURST,
       M_AWSIZE_HSIZE,
       M_AWVALID_HWRITE,
       M_BREADY,
       M_RREADY,
       M_WDATA_HWDATA,
       M_WID,
       M_WLAST,
       M_WSTRB,
       M_WVALID,
       PCIE2_LTSSM,
       PCIE2_SYSTEM_INT,
       PCIE2_WAKE_N,
       PCIE_LTSSM,
       PCIE_SYSTEM_INT,
       PLL_LOCK_INT,
       PLL_LOCKLOST_INT,
       S2_ARREADY,
       S2_AWREADY,
       S2_BID,
       S2_BRESP_HRESP,
       S2_BVALID,
       S2_RDATA_HRDATA,
       S2_RID,
       S2_RLAST,
       S2_RRESP,
       S2_RVALID,
       S2_WREADY_HREADYOUT,
       S_ARREADY,
       S_AWREADY,
       S_BID,
       S_BRESP_HRESP,
       S_BVALID,
       S_RDATA_HRDATA,
       S_RID,
       S_RLAST,
       S_RRESP,
       S_RVALID,
       S_WREADY_HREADYOUT,
       SPLL_LOCK,
       WAKE_N,
       XAUI_OUT_CLK,
       APB_CLK,
       APB_PADDR,
       APB_PENABLE,
       APB_PSEL,
       APB_PWDATA,
       APB_PWRITE,
       APB_RSTN,
       CLK_BASE,
       EPCS_PWRDN,
       EPCS_RSTN,
       EPCS_RXERR,
       EPCS_TXDATA,
       EPCS_TXOOB,
       EPCS_TXVAL,
       F2HCALIB0,
       F2HCALIB1,
       FAB_PLL_LOCK,
       FAB_REF_CLK,
       M2_ARREADY,
       M2_AWREADY,
       M2_BID,
       M2_BRESP_HRESP,
       M2_BVALID,
       M2_RDATA_HRDATA,
       M2_RID,
       M2_RLAST,
       M2_RRESP,
       M2_RVALID,
       M2_WREADY_HREADY,
       M_ARREADY,
       M_AWREADY,
       M_BID,
       M_BRESP_HRESP,
       M_BVALID,
       M_RDATA_HRDATA,
       M_RID,
       M_RLAST,
       M_RRESP,
       M_RVALID,
       M_WREADY_HREADY,
       PCIE2_INTERRUPT,
       PCIE2_PERST_N,
       PCIE2_SERDESIF_CORE_RESET_N,
       PCIE2_WAKE_REQ,
       PCIE_INTERRUPT,
       PERST_N,
       S2_ARADDR,
       S2_ARBURST,
       S2_ARID,
       S2_ARLEN,
       S2_ARLOCK,
       S2_ARSIZE,
       S2_ARVALID,
       S2_AWADDR_HADDR,
       S2_AWBURST_HTRANS,
       S2_AWID_HSEL,
       S2_AWLEN_HBURST,
       S2_AWLOCK,
       S2_AWSIZE_HSIZE,
       S2_AWVALID_HWRITE,
       S2_BREADY_HREADY,
       S2_RREADY,
       S2_WDATA_HWDATA,
       S2_WID,
       S2_WLAST,
       S2_WSTRB,
       S2_WVALID,
       S_ARADDR,
       S_ARBURST,
       S_ARID,
       S_ARLEN,
       S_ARLOCK,
       S_ARSIZE,
       S_ARVALID,
       S_AWADDR_HADDR,
       S_AWBURST_HTRANS,
       S_AWID_HSEL,
       S_AWLEN_HBURST,
       S_AWLOCK,
       S_AWSIZE_HSIZE,
       S_AWVALID_HWRITE,
       S_BREADY_HREADY,
       S_RREADY,
       S_WDATA_HWDATA,
       S_WID,
       S_WLAST,
       S_WSTRB,
       S_WVALID,
       SERDESIF_CORE_RESET_N,
       SERDESIF_PHY_RESET_N,
       WAKE_REQ,
       XAUI_FB_CLK,
       RXD3_P,
       RXD2_P,
       RXD1_P,
       RXD0_P,
       RXD3_N,
       RXD2_N,
       RXD1_N,
       RXD0_N,
       TXD3_P,
       TXD2_P,
       TXD1_P,
       TXD0_P,
       TXD3_N,
       TXD2_N,
       TXD1_N,
       TXD0_N,
       REFCLK0,
       REFCLK1
    );
output [31:0] APB_PRDATA;
output APB_PREADY;
output APB_PSLVERR;
output [1:0] ATXCLKSTABLE;
output [1:0] EPCS_READY;
output [1:0] EPCS_RXCLK;
output EPCS_RXCLK_0;
output EPCS_RXCLK_1;
output [39:0] EPCS_RXDATA;
output [1:0] EPCS_RXIDLE;
output [1:0] EPCS_RXRSTN;
output [1:0] EPCS_RXVAL;
output [1:0] EPCS_TXCLK;
output EPCS_TXCLK_0;
output EPCS_TXCLK_1;
output [1:0] EPCS_TXRSTN;
output FATC_RESET_N;
output H2FCALIB0;
output H2FCALIB1;
output [31:0] M2_ARADDR;
output [1:0] M2_ARBURST;
output [3:0] M2_ARID;
output [3:0] M2_ARLEN;
output [1:0] M2_ARSIZE;
output M2_ARVALID;
output [31:0] M2_AWADDR_HADDR;
output [1:0] M2_AWBURST_HTRANS;
output [3:0] M2_AWID;
output [3:0] M2_AWLEN_HBURST;
output [1:0] M2_AWSIZE_HSIZE;
output M2_AWVALID_HWRITE;
output M2_BREADY;
output M2_RREADY;
output [63:0] M2_WDATA_HWDATA;
output [3:0] M2_WID;
output M2_WLAST;
output [7:0] M2_WSTRB;
output M2_WVALID;
output [31:0] M_ARADDR;
output [1:0] M_ARBURST;
output [3:0] M_ARID;
output [3:0] M_ARLEN;
output [1:0] M_ARSIZE;
output M_ARVALID;
output [31:0] M_AWADDR_HADDR;
output [1:0] M_AWBURST_HTRANS;
output [3:0] M_AWID;
output [3:0] M_AWLEN_HBURST;
output [1:0] M_AWSIZE_HSIZE;
output M_AWVALID_HWRITE;
output M_BREADY;
output M_RREADY;
output [63:0] M_WDATA_HWDATA;
output [3:0] M_WID;
output M_WLAST;
output [7:0] M_WSTRB;
output M_WVALID;
output [5:0] PCIE2_LTSSM;
output PCIE2_SYSTEM_INT;
output PCIE2_WAKE_N;
output [5:0] PCIE_LTSSM;
output PCIE_SYSTEM_INT;
output PLL_LOCK_INT;
output PLL_LOCKLOST_INT;
output S2_ARREADY;
output S2_AWREADY;
output [3:0] S2_BID;
output [1:0] S2_BRESP_HRESP;
output S2_BVALID;
output [63:0] S2_RDATA_HRDATA;
output [3:0] S2_RID;
output S2_RLAST;
output [1:0] S2_RRESP;
output S2_RVALID;
output S2_WREADY_HREADYOUT;
output S_ARREADY;
output S_AWREADY;
output [3:0] S_BID;
output [1:0] S_BRESP_HRESP;
output S_BVALID;
output [63:0] S_RDATA_HRDATA;
output [3:0] S_RID;
output S_RLAST;
output [1:0] S_RRESP;
output S_RVALID;
output S_WREADY_HREADYOUT;
output SPLL_LOCK;
output WAKE_N;
output XAUI_OUT_CLK;
input  APB_CLK;
input  [14:2] APB_PADDR;
input  APB_PENABLE;
input  APB_PSEL;
input  [31:0] APB_PWDATA;
input  APB_PWRITE;
input  APB_RSTN;
input  CLK_BASE;
input  [1:0] EPCS_PWRDN;
input  [1:0] EPCS_RSTN;
input  [1:0] EPCS_RXERR;
input  [39:0] EPCS_TXDATA;
input  [1:0] EPCS_TXOOB;
input  [1:0] EPCS_TXVAL;
input  F2HCALIB0;
input  F2HCALIB1;
input  FAB_PLL_LOCK;
input  FAB_REF_CLK;
input  M2_ARREADY;
input  M2_AWREADY;
input  [3:0] M2_BID;
input  [1:0] M2_BRESP_HRESP;
input  M2_BVALID;
input  [63:0] M2_RDATA_HRDATA;
input  [3:0] M2_RID;
input  M2_RLAST;
input  [1:0] M2_RRESP;
input  M2_RVALID;
input  M2_WREADY_HREADY;
input  M_ARREADY;
input  M_AWREADY;
input  [3:0] M_BID;
input  [1:0] M_BRESP_HRESP;
input  M_BVALID;
input  [63:0] M_RDATA_HRDATA;
input  [3:0] M_RID;
input  M_RLAST;
input  [1:0] M_RRESP;
input  M_RVALID;
input  M_WREADY_HREADY;
input  [3:0] PCIE2_INTERRUPT;
input  PCIE2_PERST_N;
input  PCIE2_SERDESIF_CORE_RESET_N;
input  PCIE2_WAKE_REQ;
input  [3:0] PCIE_INTERRUPT;
input  PERST_N;
input  [31:0] S2_ARADDR;
input  [1:0] S2_ARBURST;
input  [3:0] S2_ARID;
input  [3:0] S2_ARLEN;
input  [1:0] S2_ARLOCK;
input  [1:0] S2_ARSIZE;
input  S2_ARVALID;
input  [31:0] S2_AWADDR_HADDR;
input  [1:0] S2_AWBURST_HTRANS;
input  [3:0] S2_AWID_HSEL;
input  [3:0] S2_AWLEN_HBURST;
input  [1:0] S2_AWLOCK;
input  [1:0] S2_AWSIZE_HSIZE;
input  S2_AWVALID_HWRITE;
input  S2_BREADY_HREADY;
input  S2_RREADY;
input  [63:0] S2_WDATA_HWDATA;
input  [3:0] S2_WID;
input  S2_WLAST;
input  [7:0] S2_WSTRB;
input  S2_WVALID;
input  [31:0] S_ARADDR;
input  [1:0] S_ARBURST;
input  [3:0] S_ARID;
input  [3:0] S_ARLEN;
input  [1:0] S_ARLOCK;
input  [1:0] S_ARSIZE;
input  S_ARVALID;
input  [31:0] S_AWADDR_HADDR;
input  [1:0] S_AWBURST_HTRANS;
input  [3:0] S_AWID_HSEL;
input  [3:0] S_AWLEN_HBURST;
input  [1:0] S_AWLOCK;
input  [1:0] S_AWSIZE_HSIZE;
input  S_AWVALID_HWRITE;
input  S_BREADY_HREADY;
input  S_RREADY;
input  [63:0] S_WDATA_HWDATA;
input  [3:0] S_WID;
input  S_WLAST;
input  [7:0] S_WSTRB;
input  S_WVALID;
input  SERDESIF_CORE_RESET_N;
input  SERDESIF_PHY_RESET_N;
input  WAKE_REQ;
input  XAUI_FB_CLK;
input  RXD3_P;
input  RXD2_P;
input  RXD1_P;
input  RXD0_P;
input  RXD3_N;
input  RXD2_N;
input  RXD1_N;
input  RXD0_N;
output TXD3_P;
output TXD2_P;
output TXD1_P;
output TXD0_P;
output TXD3_N;
output TXD2_N;
output TXD1_N;
output TXD0_N;
input  REFCLK0;
input  REFCLK1;

    parameter INIT = 'h0 ;
    parameter ACT_CONFIG = "" ;
    parameter ACT_SIM = 0 ;
    
endmodule


module RCOSC_25_50MHZ_FAB(
       A,
       CLKOUT
    );
input  A;
output CLKOUT;

    
endmodule


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module MSS_075(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MGPIO0B_IN,
       MGPIO10B_IN,
       MGPIO1B_IN,
       MGPIO25A_IN,
       MGPIO26A_IN,
       MGPIO27A_IN,
       MGPIO28A_IN,
       MGPIO29A_IN,
       MGPIO2B_IN,
       MGPIO30A_IN,
       MGPIO31A_IN,
       MGPIO3B_IN,
       MGPIO4B_IN,
       MGPIO5B_IN,
       MGPIO6B_IN,
       MGPIO7B_IN,
       MGPIO8B_IN,
       MGPIO9B_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_CTS_MGPIO13B_IN,
       MMUART1_DCD_MGPIO16B_IN,
       MMUART1_DSR_MGPIO14B_IN,
       MMUART1_DTR_MGPIO12B_IN,
       MMUART1_RI_MGPIO15B_IN,
       MMUART1_RTS_MGPIO11B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI0_SS4_MGPIO19A_IN,
       SPI0_SS5_MGPIO20A_IN,
       SPI0_SS6_MGPIO21A_IN,
       SPI0_SS7_MGPIO22A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       USBD_DATA0_IN,
       USBD_DATA1_IN,
       USBD_DATA2_IN,
       USBD_DATA3_IN,
       USBD_DATA4_IN,
       USBD_DATA5_IN,
       USBD_DATA6_IN,
       USBD_DATA7_MGPIO23B_IN,
       USBD_DIR_IN,
       USBD_NXT_IN,
       USBD_STP_IN,
       USBD_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MGPIO0B_OUT,
       MGPIO10B_OUT,
       MGPIO1B_OUT,
       MGPIO25A_OUT,
       MGPIO26A_OUT,
       MGPIO27A_OUT,
       MGPIO28A_OUT,
       MGPIO29A_OUT,
       MGPIO2B_OUT,
       MGPIO30A_OUT,
       MGPIO31A_OUT,
       MGPIO3B_OUT,
       MGPIO4B_OUT,
       MGPIO5B_OUT,
       MGPIO6B_OUT,
       MGPIO7B_OUT,
       MGPIO8B_OUT,
       MGPIO9B_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_CTS_MGPIO13B_OUT,
       MMUART1_DCD_MGPIO16B_OUT,
       MMUART1_DSR_MGPIO14B_OUT,
       MMUART1_DTR_MGPIO12B_OUT,
       MMUART1_RI_MGPIO15B_OUT,
       MMUART1_RTS_MGPIO11B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI0_SS4_MGPIO19A_OUT,
       SPI0_SS5_MGPIO20A_OUT,
       SPI0_SS6_MGPIO21A_OUT,
       SPI0_SS7_MGPIO22A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       USBD_DATA0_OUT,
       USBD_DATA1_OUT,
       USBD_DATA2_OUT,
       USBD_DATA3_OUT,
       USBD_DATA4_OUT,
       USBD_DATA5_OUT,
       USBD_DATA6_OUT,
       USBD_DATA7_MGPIO23B_OUT,
       USBD_DIR_OUT,
       USBD_NXT_OUT,
       USBD_STP_OUT,
       USBD_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MGPIO0B_OE,
       MGPIO10B_OE,
       MGPIO1B_OE,
       MGPIO25A_OE,
       MGPIO26A_OE,
       MGPIO27A_OE,
       MGPIO28A_OE,
       MGPIO29A_OE,
       MGPIO2B_OE,
       MGPIO30A_OE,
       MGPIO31A_OE,
       MGPIO3B_OE,
       MGPIO4B_OE,
       MGPIO5B_OE,
       MGPIO6B_OE,
       MGPIO7B_OE,
       MGPIO8B_OE,
       MGPIO9B_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_CTS_MGPIO13B_OE,
       MMUART1_DCD_MGPIO16B_OE,
       MMUART1_DSR_MGPIO14B_OE,
       MMUART1_DTR_MGPIO12B_OE,
       MMUART1_RI_MGPIO15B_OE,
       MMUART1_RTS_MGPIO11B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI0_SS4_MGPIO19A_OE,
       SPI0_SS5_MGPIO20A_OE,
       SPI0_SS6_MGPIO21A_OE,
       SPI0_SS7_MGPIO22A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE,
       USBD_DATA0_OE,
       USBD_DATA1_OE,
       USBD_DATA2_OE,
       USBD_DATA3_OE,
       USBD_DATA4_OE,
       USBD_DATA5_OE,
       USBD_DATA6_OE,
       USBD_DATA7_MGPIO23B_OE,
       USBD_DIR_OE,
       USBD_NXT_OE,
       USBD_STP_OE,
       USBD_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MGPIO0B_IN;
input  MGPIO10B_IN;
input  MGPIO1B_IN;
input  MGPIO25A_IN;
input  MGPIO26A_IN;
input  MGPIO27A_IN;
input  MGPIO28A_IN;
input  MGPIO29A_IN;
input  MGPIO2B_IN;
input  MGPIO30A_IN;
input  MGPIO31A_IN;
input  MGPIO3B_IN;
input  MGPIO4B_IN;
input  MGPIO5B_IN;
input  MGPIO6B_IN;
input  MGPIO7B_IN;
input  MGPIO8B_IN;
input  MGPIO9B_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_CTS_MGPIO13B_IN;
input  MMUART1_DCD_MGPIO16B_IN;
input  MMUART1_DSR_MGPIO14B_IN;
input  MMUART1_DTR_MGPIO12B_IN;
input  MMUART1_RI_MGPIO15B_IN;
input  MMUART1_RTS_MGPIO11B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI0_SS4_MGPIO19A_IN;
input  SPI0_SS5_MGPIO20A_IN;
input  SPI0_SS6_MGPIO21A_IN;
input  SPI0_SS7_MGPIO22A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
input  USBD_DATA0_IN;
input  USBD_DATA1_IN;
input  USBD_DATA2_IN;
input  USBD_DATA3_IN;
input  USBD_DATA4_IN;
input  USBD_DATA5_IN;
input  USBD_DATA6_IN;
input  USBD_DATA7_MGPIO23B_IN;
input  USBD_DIR_IN;
input  USBD_NXT_IN;
input  USBD_STP_IN;
input  USBD_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MGPIO0B_OUT;
output MGPIO10B_OUT;
output MGPIO1B_OUT;
output MGPIO25A_OUT;
output MGPIO26A_OUT;
output MGPIO27A_OUT;
output MGPIO28A_OUT;
output MGPIO29A_OUT;
output MGPIO2B_OUT;
output MGPIO30A_OUT;
output MGPIO31A_OUT;
output MGPIO3B_OUT;
output MGPIO4B_OUT;
output MGPIO5B_OUT;
output MGPIO6B_OUT;
output MGPIO7B_OUT;
output MGPIO8B_OUT;
output MGPIO9B_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_CTS_MGPIO13B_OUT;
output MMUART1_DCD_MGPIO16B_OUT;
output MMUART1_DSR_MGPIO14B_OUT;
output MMUART1_DTR_MGPIO12B_OUT;
output MMUART1_RI_MGPIO15B_OUT;
output MMUART1_RTS_MGPIO11B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI0_SS4_MGPIO19A_OUT;
output SPI0_SS5_MGPIO20A_OUT;
output SPI0_SS6_MGPIO21A_OUT;
output SPI0_SS7_MGPIO22A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output USBD_DATA0_OUT;
output USBD_DATA1_OUT;
output USBD_DATA2_OUT;
output USBD_DATA3_OUT;
output USBD_DATA4_OUT;
output USBD_DATA5_OUT;
output USBD_DATA6_OUT;
output USBD_DATA7_MGPIO23B_OUT;
output USBD_DIR_OUT;
output USBD_NXT_OUT;
output USBD_STP_OUT;
output USBD_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MGPIO0B_OE;
output MGPIO10B_OE;
output MGPIO1B_OE;
output MGPIO25A_OE;
output MGPIO26A_OE;
output MGPIO27A_OE;
output MGPIO28A_OE;
output MGPIO29A_OE;
output MGPIO2B_OE;
output MGPIO30A_OE;
output MGPIO31A_OE;
output MGPIO3B_OE;
output MGPIO4B_OE;
output MGPIO5B_OE;
output MGPIO6B_OE;
output MGPIO7B_OE;
output MGPIO8B_OE;
output MGPIO9B_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_CTS_MGPIO13B_OE;
output MMUART1_DCD_MGPIO16B_OE;
output MMUART1_DSR_MGPIO14B_OE;
output MMUART1_DTR_MGPIO12B_OE;
output MMUART1_RI_MGPIO15B_OE;
output MMUART1_RTS_MGPIO11B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI0_SS4_MGPIO19A_OE;
output SPI0_SS5_MGPIO20A_OE;
output SPI0_SS6_MGPIO21A_OE;
output SPI0_SS7_MGPIO22A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;
output USBD_DATA0_OE;
output USBD_DATA1_OE;
output USBD_DATA2_OE;
output USBD_DATA3_OE;
output USBD_DATA4_OE;
output USBD_DATA5_OE;
output USBD_DATA6_OE;
output USBD_DATA7_MGPIO23B_OE;
output USBD_DIR_OE;
output USBD_NXT_OE;
output USBD_STP_OE;
output USBD_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    parameter DDR_CLK_FREQ = 0.0 ;
    
endmodule


module M2S_MSS_SERDES_IF2_0_SERDES_IF2(
       M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA,
       PCIE_0_INTERRUPT_c,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR,
       APB_S_PCLK_c,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE,
       N_39,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE,
       APB_S_PRESET_N_c,
       CLK_BASE_c,
       PCIE_0_PERST_N_c,
       PCIE_0_CORE_RESET_N_c,
       PHY_RESET_N_c,
       RXD3_P,
       RXD2_P,
       RXD1_P,
       RXD0_P,
       RXD3_N,
       RXD2_N,
       RXD1_N,
       RXD0_N,
       TXD3_P,
       TXD2_P,
       TXD1_P,
       TXD0_P,
       TXD3_N,
       TXD2_N,
       TXD1_N,
       TXD0_N,
       REFCLK0_N,
       REFCLK0_P
    );
output [31:0] M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA;
input  [14:2] M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR;
input  [31:0] M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA;
input  [3:0] PCIE_0_INTERRUPT_c;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR;
input  APB_S_PCLK_c;
input  M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE;
input  N_39;
input  M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE;
input  APB_S_PRESET_N_c;
input  CLK_BASE_c;
input  PCIE_0_PERST_N_c;
input  PCIE_0_CORE_RESET_N_c;
input  PHY_RESET_N_c;
input  RXD3_P;
input  RXD2_P;
input  RXD1_P;
input  RXD0_P;
input  RXD3_N;
input  RXD2_N;
input  RXD1_N;
input  RXD0_N;
output TXD3_P;
output TXD2_P;
output TXD1_P;
output TXD0_P;
output TXD3_N;
output TXD2_N;
output TXD1_N;
output TXD0_N;
input  REFCLK0_N;
input  REFCLK0_P;

    wire VCC_net_1, GND_net_1, REFCLK0_OUT;
    
    INBUF_DIFF refclk0_inbuf_diff (.PADP(REFCLK0_P), .PADN(REFCLK0_N), 
        .Y(REFCLK0_OUT));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    SERDESIF_075 #( .INIT(1100'h080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007C0002700000000000000000000000000000000000000000000000000000007E000000000000000068400000000000000000AAB08D52278E7FF8380000000003FE1FC458F40003FFFFFBFFFFFFFFFFFFFFDFFFFFFFFFFF)
        , .ACT_CONFIG("SERDESIF_0"), .ACT_SIM(2) )  SERDESIF_INST (
        .APB_PRDATA({M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[31], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[30], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[29], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[28], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[27], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[26], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[25], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[24], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[23], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[22], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[21], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[20], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[19], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[18], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[17], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[16], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[15], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[14], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[13], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[12], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[11], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[2], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[1], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[0]}), .APB_PREADY(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY), .APB_PSLVERR(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR), .ATXCLKSTABLE({nc0, nc1})
        , .EPCS_READY({nc2, nc3}), .EPCS_RXCLK({nc4, nc5}), 
        .EPCS_RXCLK_0(), .EPCS_RXCLK_1(), .EPCS_RXDATA({nc6, nc7, nc8, 
        nc9, nc10, nc11, nc12, nc13, nc14, nc15, nc16, nc17, nc18, 
        nc19, nc20, nc21, nc22, nc23, nc24, nc25, nc26, nc27, nc28, 
        nc29, nc30, nc31, nc32, nc33, nc34, nc35, nc36, nc37, nc38, 
        nc39, nc40, nc41, nc42, nc43, nc44, nc45}), .EPCS_RXIDLE({nc46, 
        nc47}), .EPCS_RXRSTN({nc48, nc49}), .EPCS_RXVAL({nc50, nc51}), 
        .EPCS_TXCLK({nc52, nc53}), .EPCS_TXCLK_0(), .EPCS_TXCLK_1(), 
        .EPCS_TXRSTN({nc54, nc55}), .FATC_RESET_N(), .H2FCALIB0(), 
        .H2FCALIB1(), .M2_ARADDR({nc56, nc57, nc58, nc59, nc60, nc61, 
        nc62, nc63, nc64, nc65, nc66, nc67, nc68, nc69, nc70, nc71, 
        nc72, nc73, nc74, nc75, nc76, nc77, nc78, nc79, nc80, nc81, 
        nc82, nc83, nc84, nc85, nc86, nc87}), .M2_ARBURST({nc88, nc89})
        , .M2_ARID({nc90, nc91, nc92, nc93}), .M2_ARLEN({nc94, nc95, 
        nc96, nc97}), .M2_ARSIZE({nc98, nc99}), .M2_ARVALID(), 
        .M2_AWADDR_HADDR({nc100, nc101, nc102, nc103, nc104, nc105, 
        nc106, nc107, nc108, nc109, nc110, nc111, nc112, nc113, nc114, 
        nc115, nc116, nc117, nc118, nc119, nc120, nc121, nc122, nc123, 
        nc124, nc125, nc126, nc127, nc128, nc129, nc130, nc131}), 
        .M2_AWBURST_HTRANS({nc132, nc133}), .M2_AWID({nc134, nc135, 
        nc136, nc137}), .M2_AWLEN_HBURST({nc138, nc139, nc140, nc141}), 
        .M2_AWSIZE_HSIZE({nc142, nc143}), .M2_AWVALID_HWRITE(), 
        .M2_BREADY(), .M2_RREADY(), .M2_WDATA_HWDATA({nc144, nc145, 
        nc146, nc147, nc148, nc149, nc150, nc151, nc152, nc153, nc154, 
        nc155, nc156, nc157, nc158, nc159, nc160, nc161, nc162, nc163, 
        nc164, nc165, nc166, nc167, nc168, nc169, nc170, nc171, nc172, 
        nc173, nc174, nc175, nc176, nc177, nc178, nc179, nc180, nc181, 
        nc182, nc183, nc184, nc185, nc186, nc187, nc188, nc189, nc190, 
        nc191, nc192, nc193, nc194, nc195, nc196, nc197, nc198, nc199, 
        nc200, nc201, nc202, nc203, nc204, nc205, nc206, nc207}), 
        .M2_WID({nc208, nc209, nc210, nc211}), .M2_WLAST(), .M2_WSTRB({
        nc212, nc213, nc214, nc215, nc216, nc217, nc218, nc219}), 
        .M2_WVALID(), .M_ARADDR({nc220, nc221, nc222, nc223, nc224, 
        nc225, nc226, nc227, nc228, nc229, nc230, nc231, nc232, nc233, 
        nc234, nc235, nc236, nc237, nc238, nc239, nc240, nc241, nc242, 
        nc243, nc244, nc245, nc246, nc247, nc248, nc249, nc250, nc251})
        , .M_ARBURST({nc252, nc253}), .M_ARID({nc254, nc255, nc256, 
        nc257}), .M_ARLEN({nc258, nc259, nc260, nc261}), .M_ARSIZE({
        nc262, nc263}), .M_ARVALID(), .M_AWADDR_HADDR({nc264, nc265, 
        nc266, nc267, nc268, nc269, nc270, nc271, nc272, nc273, nc274, 
        nc275, nc276, nc277, nc278, nc279, nc280, nc281, nc282, nc283, 
        nc284, nc285, nc286, nc287, nc288, nc289, nc290, nc291, nc292, 
        nc293, nc294, nc295}), .M_AWBURST_HTRANS({nc296, nc297}), 
        .M_AWID({nc298, nc299, nc300, nc301}), .M_AWLEN_HBURST({nc302, 
        nc303, nc304, nc305}), .M_AWSIZE_HSIZE({nc306, nc307}), 
        .M_AWVALID_HWRITE(), .M_BREADY(), .M_RREADY(), .M_WDATA_HWDATA({
        nc308, nc309, nc310, nc311, nc312, nc313, nc314, nc315, nc316, 
        nc317, nc318, nc319, nc320, nc321, nc322, nc323, nc324, nc325, 
        nc326, nc327, nc328, nc329, nc330, nc331, nc332, nc333, nc334, 
        nc335, nc336, nc337, nc338, nc339, nc340, nc341, nc342, nc343, 
        nc344, nc345, nc346, nc347, nc348, nc349, nc350, nc351, nc352, 
        nc353, nc354, nc355, nc356, nc357, nc358, nc359, nc360, nc361, 
        nc362, nc363, nc364, nc365, nc366, nc367, nc368, nc369, nc370, 
        nc371}), .M_WID({nc372, nc373, nc374, nc375}), .M_WLAST(), 
        .M_WSTRB({nc376, nc377, nc378, nc379, nc380, nc381, nc382, 
        nc383}), .M_WVALID(), .PCIE2_LTSSM({nc384, nc385, nc386, nc387, 
        nc388, nc389}), .PCIE2_SYSTEM_INT(), .PCIE2_WAKE_N(), 
        .PCIE_LTSSM({nc390, nc391, nc392, nc393, nc394, nc395}), 
        .PCIE_SYSTEM_INT(), .PLL_LOCK_INT(), .PLL_LOCKLOST_INT(), 
        .S2_ARREADY(), .S2_AWREADY(), .S2_BID({nc396, nc397, nc398, 
        nc399}), .S2_BRESP_HRESP({nc400, nc401}), .S2_BVALID(), 
        .S2_RDATA_HRDATA({nc402, nc403, nc404, nc405, nc406, nc407, 
        nc408, nc409, nc410, nc411, nc412, nc413, nc414, nc415, nc416, 
        nc417, nc418, nc419, nc420, nc421, nc422, nc423, nc424, nc425, 
        nc426, nc427, nc428, nc429, nc430, nc431, nc432, nc433, nc434, 
        nc435, nc436, nc437, nc438, nc439, nc440, nc441, nc442, nc443, 
        nc444, nc445, nc446, nc447, nc448, nc449, nc450, nc451, nc452, 
        nc453, nc454, nc455, nc456, nc457, nc458, nc459, nc460, nc461, 
        nc462, nc463, nc464, nc465}), .S2_RID({nc466, nc467, nc468, 
        nc469}), .S2_RLAST(), .S2_RRESP({nc470, nc471}), .S2_RVALID(), 
        .S2_WREADY_HREADYOUT(), .S_ARREADY(), .S_AWREADY(), .S_BID({
        nc472, nc473, nc474, nc475}), .S_BRESP_HRESP({nc476, nc477}), 
        .S_BVALID(), .S_RDATA_HRDATA({nc478, nc479, nc480, nc481, 
        nc482, nc483, nc484, nc485, nc486, nc487, nc488, nc489, nc490, 
        nc491, nc492, nc493, nc494, nc495, nc496, nc497, nc498, nc499, 
        nc500, nc501, nc502, nc503, nc504, nc505, nc506, nc507, nc508, 
        nc509, nc510, nc511, nc512, nc513, nc514, nc515, nc516, nc517, 
        nc518, nc519, nc520, nc521, nc522, nc523, nc524, nc525, nc526, 
        nc527, nc528, nc529, nc530, nc531, nc532, nc533, nc534, nc535, 
        nc536, nc537, nc538, nc539, nc540, nc541}), .S_RID({nc542, 
        nc543, nc544, nc545}), .S_RLAST(), .S_RRESP({nc546, nc547}), 
        .S_RVALID(), .S_WREADY_HREADYOUT(), .SPLL_LOCK(), .WAKE_N(), 
        .XAUI_OUT_CLK(), .APB_CLK(APB_S_PCLK_c), .APB_PADDR({
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[14], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[13], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[12], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[11], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[2]}), .APB_PENABLE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE), .APB_PSEL(N_39), 
        .APB_PWDATA({M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[31], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[30], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[29], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[28], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[27], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[26], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[25], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[24], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[23], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[22], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[21], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[20], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[19], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[18], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[17], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[16], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[15], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[14], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[13], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[12], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[11], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[2], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[1], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[0]}), .APB_PWRITE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE), .APB_RSTN(
        APB_S_PRESET_N_c), .CLK_BASE(CLK_BASE_c), .EPCS_PWRDN({
        VCC_net_1, VCC_net_1}), .EPCS_RSTN({GND_net_1, GND_net_1}), 
        .EPCS_RXERR({VCC_net_1, VCC_net_1}), .EPCS_TXDATA({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .EPCS_TXOOB({
        VCC_net_1, VCC_net_1}), .EPCS_TXVAL({VCC_net_1, VCC_net_1}), 
        .F2HCALIB0(VCC_net_1), .F2HCALIB1(VCC_net_1), .FAB_PLL_LOCK(
        GND_net_1), .FAB_REF_CLK(VCC_net_1), .M2_ARREADY(GND_net_1), 
        .M2_AWREADY(GND_net_1), .M2_BID({VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1}), .M2_BRESP_HRESP({GND_net_1, GND_net_1})
        , .M2_BVALID(GND_net_1), .M2_RDATA_HRDATA({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .M2_RID({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .M2_RLAST(GND_net_1), 
        .M2_RRESP({GND_net_1, GND_net_1}), .M2_RVALID(GND_net_1), 
        .M2_WREADY_HREADY(GND_net_1), .M_ARREADY(GND_net_1), 
        .M_AWREADY(GND_net_1), .M_BID({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .M_BRESP_HRESP({GND_net_1, GND_net_1}), .M_BVALID(
        GND_net_1), .M_RDATA_HRDATA({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .M_RID({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .M_RLAST(GND_net_1), .M_RRESP({GND_net_1, 
        GND_net_1}), .M_RVALID(GND_net_1), .M_WREADY_HREADY(GND_net_1), 
        .PCIE2_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .PCIE2_PERST_N(GND_net_1), .PCIE2_SERDESIF_CORE_RESET_N(
        GND_net_1), .PCIE2_WAKE_REQ(VCC_net_1), .PCIE_INTERRUPT({
        PCIE_0_INTERRUPT_c[3], PCIE_0_INTERRUPT_c[2], 
        PCIE_0_INTERRUPT_c[1], PCIE_0_INTERRUPT_c[0]}), .PERST_N(
        PCIE_0_PERST_N_c), .S2_ARADDR({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .S2_ARBURST({
        GND_net_1, GND_net_1}), .S2_ARID({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .S2_ARLEN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .S2_ARLOCK({GND_net_1, GND_net_1}), 
        .S2_ARSIZE({GND_net_1, GND_net_1}), .S2_ARVALID(GND_net_1), 
        .S2_AWADDR_HADDR({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .S2_AWBURST_HTRANS({
        GND_net_1, GND_net_1}), .S2_AWID_HSEL({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .S2_AWLEN_HBURST({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .S2_AWLOCK({GND_net_1, GND_net_1}), 
        .S2_AWSIZE_HSIZE({GND_net_1, GND_net_1}), .S2_AWVALID_HWRITE(
        GND_net_1), .S2_BREADY_HREADY(GND_net_1), .S2_RREADY(GND_net_1)
        , .S2_WDATA_HWDATA({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .S2_WID({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .S2_WLAST(GND_net_1), .S2_WSTRB({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .S2_WVALID(GND_net_1), .S_ARADDR({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .S_ARBURST({GND_net_1, GND_net_1}), .S_ARID({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .S_ARLEN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .S_ARLOCK({
        GND_net_1, GND_net_1}), .S_ARSIZE({GND_net_1, GND_net_1}), 
        .S_ARVALID(GND_net_1), .S_AWADDR_HADDR({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .S_AWBURST_HTRANS({GND_net_1, GND_net_1}), .S_AWID_HSEL({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .S_AWLEN_HBURST({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .S_AWLOCK({
        GND_net_1, GND_net_1}), .S_AWSIZE_HSIZE({GND_net_1, GND_net_1})
        , .S_AWVALID_HWRITE(GND_net_1), .S_BREADY_HREADY(GND_net_1), 
        .S_RREADY(GND_net_1), .S_WDATA_HWDATA({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .S_WID({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .S_WLAST(GND_net_1), .S_WSTRB({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .S_WVALID(GND_net_1), 
        .SERDESIF_CORE_RESET_N(PCIE_0_CORE_RESET_N_c), 
        .SERDESIF_PHY_RESET_N(PHY_RESET_N_c), .WAKE_REQ(VCC_net_1), 
        .XAUI_FB_CLK(VCC_net_1), .RXD3_P(RXD3_P), .RXD2_P(RXD2_P), 
        .RXD1_P(RXD1_P), .RXD0_P(RXD0_P), .RXD3_N(RXD3_N), .RXD2_N(
        RXD2_N), .RXD1_N(RXD1_N), .RXD0_N(RXD0_N), .TXD3_P(TXD3_P), 
        .TXD2_P(TXD2_P), .TXD1_P(TXD1_P), .TXD0_P(TXD0_P), .TXD3_N(
        TXD3_N), .TXD2_N(TXD2_N), .TXD1_N(TXD1_N), .TXD0_N(TXD0_N), 
        .REFCLK0(REFCLK0_OUT), .REFCLK1(VCC_net_1));
    
endmodule


module M2S_MSS_sb_FABOSC_0_OSC(
       FABOSC_0_RCOSC_25_50MHZ_O2F,
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FABOSC_0_RCOSC_25_50MHZ_O2F;
output FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire N_RCOSC_25_50MHZ_CLKINT, GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ_FAB I_RCOSC_25_50MHZ_FAB (.A(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), .CLKOUT(
        N_RCOSC_25_50MHZ_CLKINT));
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CLKINT I_RCOSC_25_50MHZ_FAB_CLKINT (.A(N_RCOSC_25_50MHZ_CLKINT), 
        .Y(FABOSC_0_RCOSC_25_50MHZ_O2F));
    
endmodule


module CoreResetP_Z2(
       FAB_CCC_GL0_c,
       CORERESETP_0_SDIF_RELEASED,
       FABOSC_0_RCOSC_25_50MHZ_O2F,
       INIT_DONE_int,
       SYSRESET_POR,
       M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F,
       MSS_ADLIB_INST_RNI7K43,
       CORECONFIGP_0_CONFIG1_DONE,
       CORECONFIGP_0_CONFIG2_DONE,
       SDIF0_SPLL_LOCK_c,
       CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET,
       SDIF0_1_CORE_RESET_N_c,
       CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET,
       SDIF0_0_CORE_RESET_N_c,
       CORECONFIGP_0_SOFT_SDIF0_PHY_RESET,
       SDIF0_PHY_RESET_N_c
    );
input  FAB_CCC_GL0_c;
output CORERESETP_0_SDIF_RELEASED;
input  FABOSC_0_RCOSC_25_50MHZ_O2F;
output INIT_DONE_int;
input  SYSRESET_POR;
input  M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F;
input  MSS_ADLIB_INST_RNI7K43;
input  CORECONFIGP_0_CONFIG1_DONE;
input  CORECONFIGP_0_CONFIG2_DONE;
input  SDIF0_SPLL_LOCK_c;
input  CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET;
output SDIF0_1_CORE_RESET_N_c;
input  CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET;
output SDIF0_0_CORE_RESET_N_c;
input  CORECONFIGP_0_SOFT_SDIF0_PHY_RESET;
output SDIF0_PHY_RESET_N_c;

    wire sm0_areset_n_clk_base, sdif0_areset_n_clk_base_net_1, 
        sm0_areset_n_rcosc, sdif0_areset_n_rcosc_net_1, 
        \count_sdif0[0]_net_1 , \count_sdif0_s[0] , 
        \count_ddr[0]_net_1 , \count_ddr_s[0] , \sdif0_state[0]_net_1 , 
        \sdif0_state_i_0[0] , count_sdif0_enable_net_1, VCC_net_1, 
        N_11, GND_net_1, next_sdif_released_0_sqmuxa, 
        ddr_settled_net_1, ddr_settled4_net_1, 
        release_sdif0_core_net_1, release_sdif0_core4_net_1, 
        SDIF0_PHY_RESET_N_int_net_1, next_sdif0_phy_reset_n_0_sqmuxa, 
        SDIF0_CORE_RESET_N_0_net_1, N_28, count_ddr_enable_net_1, 
        next_count_ddr_enable_0_sqmuxa, 
        un1_next_ddr_ready_0_sqmuxa_0_net_1, mss_ready_select_net_1, 
        POWER_ON_RESET_N_clk_base_net_1, mss_ready_select4_net_1, 
        \sm0_state[6]_net_1 , mss_ready_state_net_1, 
        RESET_N_M2F_clk_base_net_1, N_8, \sdif0_state[1]_net_1 , 
        N_4_i_0, \sm0_state[3]_net_1 , \sm0_state_ns[3] , 
        \sm0_state[4]_net_1 , \sm0_state_ns[4] , \sm0_state[5]_net_1 , 
        \sm0_state_ns[5] , N_19_i_0, \sm0_state[0]_net_1 , 
        \sm0_state[1]_net_1 , \sm0_state[2]_net_1 , 
        \sm0_state_ns[2]_net_1 , release_sdif3_core_clk_base, 
        release_sdif3_core_q1, POWER_ON_RESET_N_q1_net_1, 
        RESET_N_M2F_q1_net_1, FIC_2_APB_M_PRESET_N_clk_base_net_1, 
        FIC_2_APB_M_PRESET_N_q1_net_1, sm0_areset_n_q1_net_1, 
        sm0_areset_n_i_0_i, sm0_areset_n_rcosc_q1_net_1, 
        MSS_HPMS_READY_int_net_1, MSS_HPMS_READY_int_4_net_1, 
        count_ddr_enable_q1_net_1, count_sdif0_enable_q1_net_1, 
        ddr_settled_q1_net_1, release_sdif0_core_q1_net_1, 
        release_sdif2_core, sdif3_spll_lock_q1_net_1, 
        sdif0_spll_lock_q2_net_1, sdif0_spll_lock_q1_net_1, 
        count_ddr_enable_rcosc_net_1, count_sdif0_enable_rcosc_net_1, 
        ddr_settled_clk_base_net_1, release_sdif0_core_clk_base_net_1, 
        CONFIG1_DONE_clk_base_net_1, CONFIG1_DONE_q1_net_1, 
        CONFIG2_DONE_clk_base_net_1, CONFIG2_DONE_q1_net_1, 
        sdif3_spll_lock_q2_net_1, \count_ddr[1]_net_1 , 
        \count_ddr_s[1] , \count_ddr[2]_net_1 , \count_ddr_s[2] , 
        \count_ddr[3]_net_1 , \count_ddr_s[3] , \count_ddr[4]_net_1 , 
        \count_ddr_s[4] , \count_ddr[5]_net_1 , \count_ddr_s[5] , 
        \count_ddr[6]_net_1 , \count_ddr_s[6] , \count_ddr[7]_net_1 , 
        \count_ddr_s[7] , \count_ddr[8]_net_1 , \count_ddr_s[8] , 
        \count_ddr[9]_net_1 , \count_ddr_s[9] , \count_ddr[10]_net_1 , 
        \count_ddr_s[10] , \count_ddr[11]_net_1 , \count_ddr_s[11] , 
        \count_ddr[12]_net_1 , \count_ddr_s[12] , 
        \count_ddr[13]_net_1 , \count_ddr_s[13]_net_1 , 
        \count_sdif0[1]_net_1 , \count_sdif0_s[1] , 
        \count_sdif0[2]_net_1 , \count_sdif0_s[2] , 
        \count_sdif0[3]_net_1 , \count_sdif0_s[3] , 
        \count_sdif0[4]_net_1 , \count_sdif0_s[4] , 
        \count_sdif0[5]_net_1 , \count_sdif0_s[5] , 
        \count_sdif0[6]_net_1 , \count_sdif0_s[6] , 
        \count_sdif0[7]_net_1 , \count_sdif0_s[7] , 
        \count_sdif0[8]_net_1 , \count_sdif0_s[8] , 
        \count_sdif0[9]_net_1 , \count_sdif0_s[9] , 
        \count_sdif0[10]_net_1 , \count_sdif0_s[10] , 
        \count_sdif0[11]_net_1 , \count_sdif0_s[11] , 
        \count_sdif0[12]_net_1 , \count_sdif0_s[12]_net_1 , 
        count_sdif0_s_142_FCO, \count_sdif0_cry[1]_net_1 , 
        \count_sdif0_cry[2]_net_1 , \count_sdif0_cry[3]_net_1 , 
        \count_sdif0_cry[4]_net_1 , \count_sdif0_cry[5]_net_1 , 
        \count_sdif0_cry[6]_net_1 , \count_sdif0_cry[7]_net_1 , 
        \count_sdif0_cry[8]_net_1 , \count_sdif0_cry[9]_net_1 , 
        \count_sdif0_cry[10]_net_1 , \count_sdif0_cry[11]_net_1 , 
        count_ddr_s_143_FCO, \count_ddr_cry[1]_net_1 , 
        \count_ddr_cry[2]_net_1 , \count_ddr_cry[3]_net_1 , 
        \count_ddr_cry[4]_net_1 , \count_ddr_cry[5]_net_1 , 
        \count_ddr_cry[6]_net_1 , \count_ddr_cry[7]_net_1 , 
        \count_ddr_cry[8]_net_1 , \count_ddr_cry[9]_net_1 , 
        \count_ddr_cry[10]_net_1 , \count_ddr_cry[11]_net_1 , 
        \count_ddr_cry[12]_net_1 , release_sdif0_core4_1_net_1, 
        release_sdif0_core4_7_net_1, release_sdif0_core4_8_net_1, 
        ddr_settled4_6_net_1, N_25, ddr_settled4_9_net_1, 
        ddr_settled4_8_net_1, ddr_settled4_7_net_1, N_26;
    
    SLE \sdif0_state[0]  (.D(N_8), .CLK(FAB_CCC_GL0_c), .EN(VCC_net_1), 
        .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\sdif0_state[0]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \sm0_state_ns_0_o2[3]  (.A(
        sdif0_spll_lock_q2_net_1), .B(sdif3_spll_lock_q2_net_1), .Y(
        N_25));
    CFG1 #( .INIT(2'h1) )  count_sdif0_enable_RNO (.A(
        \sdif0_state[0]_net_1 ), .Y(\sdif0_state_i_0[0] ));
    SLE sdif3_spll_lock_q2 (.D(sdif3_spll_lock_q1_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(sdif3_spll_lock_q2_net_1));
    SLE \count_ddr[5]  (.D(\count_ddr_s[5] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[5]_net_1 ));
    SLE count_sdif0_enable_q1 (.D(count_sdif0_enable_net_1), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(VCC_net_1), .ALn(
        sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(count_sdif0_enable_q1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[2]  (.A(VCC_net_1), .B(
        \count_ddr[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[1]_net_1 ), .S(\count_ddr_s[2] ), .Y(), .FCO(
        \count_ddr_cry[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  MSS_HPMS_READY_int_RNITK3D (.A(SYSRESET_POR)
        , .B(MSS_HPMS_READY_int_net_1), .Y(sm0_areset_n_i_0_i));
    CFG4 #( .INIT(16'h0001) )  ddr_settled4_8 (.A(
        \count_ddr[12]_net_1 ), .B(\count_ddr[7]_net_1 ), .C(
        \count_ddr[5]_net_1 ), .D(\count_ddr[1]_net_1 ), .Y(
        ddr_settled4_8_net_1));
    SLE \count_sdif0[8]  (.D(\count_sdif0_s[8] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[8]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[1]  (.A(VCC_net_1), .B(
        \count_ddr[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        count_ddr_s_143_FCO), .S(\count_ddr_s[1] ), .Y(), .FCO(
        \count_ddr_cry[1]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  release_sdif0_core4 (.A(
        release_sdif0_core4_1_net_1), .B(release_sdif0_core4_7_net_1), 
        .C(\count_sdif0[6]_net_1 ), .D(release_sdif0_core4_8_net_1), 
        .Y(release_sdif0_core4_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_s[13]  (.A(VCC_net_1), .B(
        \count_ddr[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[12]_net_1 ), .S(\count_ddr_s[13]_net_1 ), .Y(), 
        .FCO());
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[1]  (.A(VCC_net_1), 
        .B(\count_sdif0[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        count_sdif0_s_142_FCO), .S(\count_sdif0_s[1] ), .Y(), .FCO(
        \count_sdif0_cry[1]_net_1 ));
    SLE POWER_ON_RESET_N_q1 (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        VCC_net_1), .ALn(SYSRESET_POR), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_q1_net_1));
    SLE \count_ddr[13]  (.D(\count_ddr_s[13]_net_1 ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[13]_net_1 ));
    SLE \count_ddr[12]  (.D(\count_ddr_s[12] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[12]_net_1 ));
    CFG4 #( .INIT(16'h7FFF) )  release_sdif0_core4_1 (.A(
        \count_sdif0[11]_net_1 ), .B(\count_sdif0[8]_net_1 ), .C(
        \count_sdif0[5]_net_1 ), .D(\count_sdif0[2]_net_1 ), .Y(
        release_sdif0_core4_1_net_1));
    SLE SDIF0_CORE_RESET_N_0 (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        N_28), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        SDIF0_CORE_RESET_N_0_net_1));
    SLE \sm0_state[6]  (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        N_19_i_0), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sm0_state[6]_net_1 ));
    SLE \sm0_state[4]  (.D(\sm0_state_ns[4] ), .CLK(FAB_CCC_GL0_c), 
        .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sm0_state[4]_net_1 ));
    CFG3 #( .INIT(8'hE0) )  MSS_HPMS_READY_int_4 (.A(
        RESET_N_M2F_clk_base_net_1), .B(mss_ready_select_net_1), .C(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .Y(
        MSS_HPMS_READY_int_4_net_1));
    SLE ddr_settled (.D(VCC_net_1), .CLK(FABOSC_0_RCOSC_25_50MHZ_O2F), 
        .EN(ddr_settled4_net_1), .ALn(sm0_areset_n_rcosc), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(ddr_settled_net_1));
    SLE sdif0_areset_n_rcosc (.D(sm0_areset_n_rcosc_q1_net_1), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(VCC_net_1), .ALn(
        sm0_areset_n_i_0_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(sdif0_areset_n_rcosc_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[6]  (.A(VCC_net_1), 
        .B(\count_sdif0[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[5]_net_1 ), .S(\count_sdif0_s[6] ), .Y(), 
        .FCO(\count_sdif0_cry[6]_net_1 ));
    CFG2 #( .INIT(4'h4) )  SDIF0_PHY_RESET_N (.A(
        CORECONFIGP_0_SOFT_SDIF0_PHY_RESET), .B(
        SDIF0_PHY_RESET_N_int_net_1), .Y(SDIF0_PHY_RESET_N_c));
    GND GND (.Y(GND_net_1));
    SLE sdif0_areset_n_clk_base (.D(sm0_areset_n_q1_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_i_0_i), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(sdif0_areset_n_clk_base_net_1));
    CFG1 #( .INIT(2'h1) )  \count_ddr_RNO[0]  (.A(\count_ddr[0]_net_1 )
        , .Y(\count_ddr_s[0] ));
    SLE \count_ddr[11]  (.D(\count_ddr_s[11] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[11]_net_1 ));
    SLE ddr_settled_clk_base (.D(ddr_settled_q1_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(ddr_settled_clk_base_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[9]  (.A(VCC_net_1), 
        .B(\count_sdif0[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[8]_net_1 ), .S(\count_sdif0_s[9] ), .Y(), 
        .FCO(\count_sdif0_cry[9]_net_1 ));
    SLE release_sdif0_core_q1 (.D(release_sdif0_core_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(release_sdif0_core_q1_net_1));
    SLE \sm0_state[0]  (.D(GND_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sm0_state[0]_net_1 ));
    CLKINT sdif0_areset_n_clk_base_RNI7MR6 (.A(
        sdif0_areset_n_clk_base_net_1), .Y(sm0_areset_n_clk_base));
    SLE \sm0_state[3]  (.D(\sm0_state_ns[3] ), .CLK(FAB_CCC_GL0_c), 
        .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sm0_state[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[4]  (.A(VCC_net_1), 
        .B(\count_sdif0[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[3]_net_1 ), .S(\count_sdif0_s[4] ), .Y(), 
        .FCO(\count_sdif0_cry[4]_net_1 ));
    SLE \sm0_state[5]  (.D(\sm0_state_ns[5] ), .CLK(FAB_CCC_GL0_c), 
        .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sm0_state[5]_net_1 ));
    SLE \count_sdif0[2]  (.D(\count_sdif0_s[2] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[2]_net_1 ));
    SLE \count_ddr[10]  (.D(\count_ddr_s[10] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[10]_net_1 ));
    SLE \count_ddr[7]  (.D(\count_ddr_s[7] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[7]_net_1 ));
    SLE INIT_DONE_int_inst_1 (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        \sm0_state[6]_net_1 ), .ALn(sm0_areset_n_clk_base), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(INIT_DONE_int));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[9]  (.A(VCC_net_1), .B(
        \count_ddr[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[8]_net_1 ), .S(\count_ddr_s[9] ), .Y(), .FCO(
        \count_ddr_cry[9]_net_1 ));
    SLE SDIF_RELEASED_int (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        next_sdif_released_0_sqmuxa), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CORERESETP_0_SDIF_RELEASED));
    CFG4 #( .INIT(16'hECA0) )  un1_next_ddr_ready_0_sqmuxa_0 (.A(
        \sm0_state[3]_net_1 ), .B(ddr_settled_clk_base_net_1), .C(
        sdif3_spll_lock_q2_net_1), .D(\sm0_state[4]_net_1 ), .Y(
        un1_next_ddr_ready_0_sqmuxa_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[10]  (.A(VCC_net_1), 
        .B(\count_sdif0[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\count_sdif0_cry[9]_net_1 ), .S(\count_sdif0_s[10] ), .Y()
        , .FCO(\count_sdif0_cry[10]_net_1 ));
    CFG4 #( .INIT(16'hC0EA) )  \sm0_state_ns_0[4]  (.A(
        \sm0_state[3]_net_1 ), .B(\sm0_state[4]_net_1 ), .C(N_26), .D(
        N_25), .Y(\sm0_state_ns[4] ));
    VCC VCC (.Y(VCC_net_1));
    SLE sm0_areset_n_q1 (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        VCC_net_1), .ALn(sm0_areset_n_i_0_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sm0_areset_n_q1_net_1));
    SLE sdif0_spll_lock_q1 (.D(SDIF0_SPLL_LOCK_c), .CLK(FAB_CCC_GL0_c), 
        .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sdif0_spll_lock_q1_net_1));
    SLE release_sdif0_core (.D(VCC_net_1), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(release_sdif0_core4_net_1), 
        .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(release_sdif0_core_net_1));
    SLE \count_sdif0[11]  (.D(\count_sdif0_s[11] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[11]_net_1 ));
    SLE MSS_HPMS_READY_int (.D(MSS_HPMS_READY_int_4_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        MSS_HPMS_READY_int_net_1));
    SLE SDIF0_PHY_RESET_N_int (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        next_sdif0_phy_reset_n_0_sqmuxa), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(SDIF0_PHY_RESET_N_int_net_1));
    CFG4 #( .INIT(16'h8000) )  \sm0_state_ns_0_a2_0[5]  (.A(
        \sm0_state[4]_net_1 ), .B(ddr_settled_clk_base_net_1), .C(
        release_sdif3_core_clk_base), .D(
        release_sdif0_core_clk_base_net_1), .Y(
        next_sdif_released_0_sqmuxa));
    CFG2 #( .INIT(4'h4) )  SDIF0_1_CORE_RESET_N_0_a2 (.A(
        CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET), .B(
        SDIF0_CORE_RESET_N_0_net_1), .Y(SDIF0_1_CORE_RESET_N_c));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[2]  (.A(VCC_net_1), 
        .B(\count_sdif0[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[1]_net_1 ), .S(\count_sdif0_s[2] ), .Y(), 
        .FCO(\count_sdif0_cry[2]_net_1 ));
    SLE CONFIG2_DONE_q1 (.D(CORECONFIGP_0_CONFIG2_DONE), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CONFIG2_DONE_q1_net_1));
    CFG3 #( .INIT(8'hF2) )  \sm0_state_ns[2]  (.A(\sm0_state[2]_net_1 )
        , .B(CONFIG1_DONE_clk_base_net_1), .C(\sm0_state[1]_net_1 ), 
        .Y(\sm0_state_ns[2]_net_1 ));
    SLE \count_ddr[0]  (.D(\count_ddr_s[0] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[0]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \sm0_state_ns_0[3]  (.A(
        CONFIG1_DONE_clk_base_net_1), .B(N_25), .C(
        \sm0_state[2]_net_1 ), .D(\sm0_state[3]_net_1 ), .Y(
        \sm0_state_ns[3] ));
    CFG4 #( .INIT(16'h8000) )  next_sdif0_core_reset_n_0_sqmuxa_i_i_a2 
        (.A(release_sdif0_core_clk_base_net_1), .B(
        \sdif0_state[1]_net_1 ), .C(ddr_settled_clk_base_net_1), .D(
        \sdif0_state[0]_net_1 ), .Y(N_28));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[4]  (.A(VCC_net_1), .B(
        \count_ddr[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[3]_net_1 ), .S(\count_ddr_s[4] ), .Y(), .FCO(
        \count_ddr_cry[4]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  release_sdif0_core4_7 (.A(
        \count_sdif0[10]_net_1 ), .B(\count_sdif0[9]_net_1 ), .C(
        \count_sdif0[7]_net_1 ), .D(\count_sdif0[0]_net_1 ), .Y(
        release_sdif0_core4_7_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[5]  (.A(VCC_net_1), 
        .B(\count_sdif0[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[4]_net_1 ), .S(\count_sdif0_s[5] ), .Y(), 
        .FCO(\count_sdif0_cry[5]_net_1 ));
    SLE sdif0_spll_lock_q2 (.D(sdif0_spll_lock_q1_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(sdif0_spll_lock_q2_net_1));
    SLE \count_ddr[2]  (.D(\count_ddr_s[2] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[2]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  count_sdif0_s_142 (.A(VCC_net_1), .B(
        \count_sdif0[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(count_sdif0_s_142_FCO));
    SLE RESET_N_M2F_q1 (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        VCC_net_1), .ALn(M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(RESET_N_M2F_q1_net_1));
    SLE count_sdif0_enable_rcosc (.D(count_sdif0_enable_q1_net_1), 
        .CLK(FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(VCC_net_1), .ALn(
        sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(count_sdif0_enable_rcosc_net_1)
        );
    SLE \sm0_state[2]  (.D(\sm0_state_ns[2]_net_1 ), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\sm0_state[2]_net_1 ));
    SLE \sm0_state[1]  (.D(\sm0_state[0]_net_1 ), .CLK(FAB_CCC_GL0_c), 
        .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sm0_state[1]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  release_sdif0_core4_8 (.A(
        \count_sdif0[12]_net_1 ), .B(\count_sdif0[4]_net_1 ), .C(
        \count_sdif0[3]_net_1 ), .D(\count_sdif0[1]_net_1 ), .Y(
        release_sdif0_core4_8_net_1));
    SLE count_ddr_enable_q1 (.D(count_ddr_enable_net_1), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(VCC_net_1), .ALn(
        sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(count_ddr_enable_q1_net_1));
    SLE release_sdif1_core_clk_base (.D(release_sdif3_core_q1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(release_sdif3_core_clk_base));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[7]  (.A(VCC_net_1), .B(
        \count_ddr[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[6]_net_1 ), .S(\count_ddr_s[7] ), .Y(), .FCO(
        \count_ddr_cry[7]_net_1 ));
    SLE CONFIG1_DONE_q1 (.D(CORECONFIGP_0_CONFIG1_DONE), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CONFIG1_DONE_q1_net_1));
    SLE \count_ddr[6]  (.D(\count_ddr_s[6] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[6]_net_1 ));
    SLE count_ddr_enable_rcosc (.D(count_ddr_enable_q1_net_1), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(VCC_net_1), .ALn(
        sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(count_ddr_enable_rcosc_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[12]  (.A(VCC_net_1), .B(
        \count_ddr[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[11]_net_1 ), .S(\count_ddr_s[12] ), .Y(), .FCO(
        \count_ddr_cry[12]_net_1 ));
    CFG2 #( .INIT(4'hE) )  un1_next_sdif0_core_reset_n_0_sqmuxa_i_i (
        .A(next_sdif0_phy_reset_n_0_sqmuxa), .B(N_28), .Y(N_11));
    CFG4 #( .INIT(16'h0001) )  ddr_settled4_9 (.A(\count_ddr[6]_net_1 )
        , .B(\count_ddr[3]_net_1 ), .C(\count_ddr[2]_net_1 ), .D(
        \count_ddr[0]_net_1 ), .Y(ddr_settled4_9_net_1));
    SLE \count_sdif0[1]  (.D(\count_sdif0_s[1] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[1]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[6]  (.A(VCC_net_1), .B(
        \count_ddr[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[5]_net_1 ), .S(\count_ddr_s[6] ), .Y(), .FCO(
        \count_ddr_cry[6]_net_1 ));
    SLE ddr_settled_q1 (.D(ddr_settled_net_1), .CLK(FAB_CCC_GL0_c), 
        .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        ddr_settled_q1_net_1));
    CFG2 #( .INIT(4'h4) )  SDIF0_0_CORE_RESET_N_0_a2 (.A(
        CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET), .B(
        SDIF0_CORE_RESET_N_0_net_1), .Y(SDIF0_0_CORE_RESET_N_c));
    SLE \count_sdif0[4]  (.D(\count_sdif0_s[4] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[4]_net_1 ));
    SLE \count_sdif0[5]  (.D(\count_sdif0_s[5] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[5]_net_1 ));
    CFG2 #( .INIT(4'h8) )  mss_ready_select4 (.A(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .B(mss_ready_state_net_1)
        , .Y(mss_ready_select4_net_1));
    SLE FIC_2_APB_M_PRESET_N_q1 (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), 
        .EN(VCC_net_1), .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        FIC_2_APB_M_PRESET_N_q1_net_1));
    SLE \count_sdif0[10]  (.D(\count_sdif0_s[10] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[10]_net_1 ));
    SLE CONFIG1_DONE_clk_base (.D(CONFIG1_DONE_q1_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CONFIG1_DONE_clk_base_net_1));
    SLE \count_ddr[8]  (.D(\count_ddr_s[8] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[8]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[3]  (.A(VCC_net_1), .B(
        \count_ddr[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[2]_net_1 ), .S(\count_ddr_s[3] ), .Y(), .FCO(
        \count_ddr_cry[3]_net_1 ));
    SLE release_sdif1_core (.D(VCC_net_1), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(VCC_net_1), .ALn(
        sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(release_sdif2_core));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_s[12]  (.A(VCC_net_1), .B(
        \count_sdif0[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[11]_net_1 ), .S(\count_sdif0_s[12]_net_1 ), 
        .Y(), .FCO());
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[11]  (.A(VCC_net_1), .B(
        \count_ddr[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[10]_net_1 ), .S(\count_ddr_s[11] ), .Y(), .FCO(
        \count_ddr_cry[11]_net_1 ));
    SLE CONFIG2_DONE_clk_base (.D(CONFIG2_DONE_q1_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(CONFIG2_DONE_clk_base_net_1));
    SLE \count_sdif0[0]  (.D(\count_sdif0_s[0] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[0]_net_1 ));
    SLE \count_sdif0[12]  (.D(\count_sdif0_s[12]_net_1 ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[12]_net_1 ));
    SLE \count_ddr[3]  (.D(\count_ddr_s[3] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[3]_net_1 ));
    SLE release_sdif1_core_q1 (.D(release_sdif2_core), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(sm0_areset_n_clk_base), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(release_sdif3_core_q1));
    SLE \count_ddr[4]  (.D(\count_ddr_s[4] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[4]_net_1 ));
    SLE mss_ready_select (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        mss_ready_select4_net_1), .ALn(POWER_ON_RESET_N_clk_base_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(mss_ready_select_net_1));
    CFG4 #( .INIT(16'hCCB3) )  \sdif0_state_ns_1_0_.m2_i  (.A(
        sdif0_spll_lock_q2_net_1), .B(\sdif0_state[1]_net_1 ), .C(
        CONFIG1_DONE_clk_base_net_1), .D(\sdif0_state[0]_net_1 ), .Y(
        N_8));
    SLE \count_sdif0[7]  (.D(\count_sdif0_s[7] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[7]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  count_ddr_s_143 (.A(VCC_net_1), .B(
        \count_ddr[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(count_ddr_s_143_FCO));
    SLE POWER_ON_RESET_N_clk_base (.D(POWER_ON_RESET_N_q1_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(SYSRESET_POR), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(POWER_ON_RESET_N_clk_base_net_1));
    CFG4 #( .INIT(16'h0080) )  
        un1_next_sdif0_core_reset_n_0_sqmuxa_i_i_a2 (.A(
        sdif0_spll_lock_q2_net_1), .B(\sdif0_state[1]_net_1 ), .C(
        CONFIG1_DONE_clk_base_net_1), .D(\sdif0_state[0]_net_1 ), .Y(
        next_sdif0_phy_reset_n_0_sqmuxa));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[5]  (.A(VCC_net_1), .B(
        \count_ddr[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[4]_net_1 ), .S(\count_ddr_s[5] ), .Y(), .FCO(
        \count_ddr_cry[5]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \sdif0_state_ns_1_0_.N_4_i  (.A(
        \sdif0_state[0]_net_1 ), .B(\sdif0_state[1]_net_1 ), .Y(
        N_4_i_0));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[11]  (.A(VCC_net_1), 
        .B(\count_sdif0[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(\count_sdif0_cry[10]_net_1 ), .S(\count_sdif0_s[11] ), .Y(
        ), .FCO(\count_sdif0_cry[11]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[7]  (.A(VCC_net_1), 
        .B(\count_sdif0[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[6]_net_1 ), .S(\count_sdif0_s[7] ), .Y(), 
        .FCO(\count_sdif0_cry[7]_net_1 ));
    SLE \count_ddr[9]  (.D(\count_ddr_s[9] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[9]_net_1 ));
    SLE \sdif0_state[1]  (.D(N_4_i_0), .CLK(FAB_CCC_GL0_c), .EN(
        VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \sdif0_state[1]_net_1 ));
    SLE sm0_areset_n_rcosc_q1 (.D(VCC_net_1), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(VCC_net_1), .ALn(
        sm0_areset_n_i_0_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(sm0_areset_n_rcosc_q1_net_1));
    CFG2 #( .INIT(4'h8) )  \sm0_state_RNO[6]  (.A(
        CONFIG2_DONE_clk_base_net_1), .B(\sm0_state[5]_net_1 ), .Y(
        N_19_i_0));
    CFG2 #( .INIT(4'h4) )  ddr_settled4_6 (.A(\count_ddr[11]_net_1 ), 
        .B(\count_ddr[13]_net_1 ), .Y(ddr_settled4_6_net_1));
    SLE count_ddr_enable (.D(next_count_ddr_enable_0_sqmuxa), .CLK(
        FAB_CCC_GL0_c), .EN(un1_next_ddr_ready_0_sqmuxa_0_net_1), .ALn(
        sm0_areset_n_clk_base), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(count_ddr_enable_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[8]  (.A(VCC_net_1), 
        .B(\count_sdif0[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[7]_net_1 ), .S(\count_sdif0_s[8] ), .Y(), 
        .FCO(\count_sdif0_cry[8]_net_1 ));
    SLE \count_sdif0[6]  (.D(\count_sdif0_s[6] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[6]_net_1 ));
    SLE \count_sdif0[9]  (.D(\count_sdif0_s[9] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[9]_net_1 ));
    SLE release_sdif0_core_clk_base (.D(release_sdif0_core_q1_net_1), 
        .CLK(FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(
        sm0_areset_n_clk_base), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        release_sdif0_core_clk_base_net_1));
    CFG1 #( .INIT(2'h1) )  \count_sdif0_RNO[0]  (.A(
        \count_sdif0[0]_net_1 ), .Y(\count_sdif0_s[0] ));
    SLE \count_sdif0[3]  (.D(\count_sdif0_s[3] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(
        count_sdif0_enable_rcosc_net_1), .ALn(sm0_areset_n_rcosc), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\count_sdif0[3]_net_1 ));
    CLKINT sdif0_areset_n_rcosc_RNIDB37 (.A(sdif0_areset_n_rcosc_net_1)
        , .Y(sm0_areset_n_rcosc));
    CFG2 #( .INIT(4'h8) )  un1_next_ddr_ready_0_sqmuxa_0_a2_0 (.A(
        \sm0_state[3]_net_1 ), .B(sdif3_spll_lock_q2_net_1), .Y(
        next_count_ddr_enable_0_sqmuxa));
    SLE RESET_N_M2F_clk_base (.D(RESET_N_M2F_q1_net_1), .CLK(
        FAB_CCC_GL0_c), .EN(VCC_net_1), .ALn(
        M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RESET_N_M2F_clk_base_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[10]  (.A(VCC_net_1), .B(
        \count_ddr[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[9]_net_1 ), .S(\count_ddr_s[10] ), .Y(), .FCO(
        \count_ddr_cry[10]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  ddr_settled4_7 (.A(
        \count_ddr[10]_net_1 ), .B(\count_ddr[9]_net_1 ), .C(
        \count_ddr[8]_net_1 ), .D(\count_ddr[4]_net_1 ), .Y(
        ddr_settled4_7_net_1));
    SLE count_sdif0_enable (.D(\sdif0_state_i_0[0] ), .CLK(
        FAB_CCC_GL0_c), .EN(N_11), .ALn(sm0_areset_n_clk_base), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(count_sdif0_enable_net_1));
    CFG4 #( .INIT(16'h8000) )  ddr_settled4 (.A(ddr_settled4_6_net_1), 
        .B(ddr_settled4_7_net_1), .C(ddr_settled4_8_net_1), .D(
        ddr_settled4_9_net_1), .Y(ddr_settled4_net_1));
    SLE sdif3_spll_lock_q1 (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        VCC_net_1), .ALn(sm0_areset_n_clk_base), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        sdif3_spll_lock_q1_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_sdif0_cry[3]  (.A(VCC_net_1), 
        .B(\count_sdif0[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_sdif0_cry[2]_net_1 ), .S(\count_sdif0_s[3] ), .Y(), 
        .FCO(\count_sdif0_cry[3]_net_1 ));
    CFG3 #( .INIT(8'hAE) )  \sm0_state_ns_0[5]  (.A(
        next_sdif_released_0_sqmuxa), .B(\sm0_state[5]_net_1 ), .C(
        CONFIG2_DONE_clk_base_net_1), .Y(\sm0_state_ns[5] ));
    SLE FIC_2_APB_M_PRESET_N_clk_base (.D(
        FIC_2_APB_M_PRESET_N_q1_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        VCC_net_1), .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        FIC_2_APB_M_PRESET_N_clk_base_net_1));
    SLE mss_ready_state (.D(VCC_net_1), .CLK(FAB_CCC_GL0_c), .EN(
        RESET_N_M2F_clk_base_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        mss_ready_state_net_1));
    ARI1 #( .INIT(20'h4AA00) )  \count_ddr_cry[8]  (.A(VCC_net_1), .B(
        \count_ddr[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        \count_ddr_cry[7]_net_1 ), .S(\count_ddr_s[8] ), .Y(), .FCO(
        \count_ddr_cry[8]_net_1 ));
    SLE \count_ddr[1]  (.D(\count_ddr_s[1] ), .CLK(
        FABOSC_0_RCOSC_25_50MHZ_O2F), .EN(count_ddr_enable_rcosc_net_1)
        , .ALn(sm0_areset_n_rcosc), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\count_ddr[1]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \sm0_state_ns_0_o2[4]  (.A(
        release_sdif3_core_clk_base), .B(
        release_sdif0_core_clk_base_net_1), .C(
        ddr_settled_clk_base_net_1), .Y(N_26));
    
endmodule


module M2S_MSS_sb_MSS(
       MDDR_DQ,
       MDDR_DM_RDQS,
       MDDR_BA,
       MDDR_ADDR,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA,
       CORECONFIGP_0_MDDR_APBmslave_PRDATA,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA,
       MDDR_DQS_N,
       MDDR_DQS,
       FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA,
       MSS_ADLIB_INST_RNI7K43,
       un1_M2S_MSS_sb_0_4_i_0,
       SPI_1_SS0,
       SPI_1_DO,
       SPI_1_DI,
       SPI_1_CLK,
       SPI_0_SS0,
       SPI_0_DO,
       SPI_0_DI,
       SPI_0_CLK,
       MMUART_1_TXD,
       MMUART_1_RXD,
       MMUART_0_TXD,
       MMUART_0_RXD,
       MDDR_WE_N,
       MDDR_RESET_N,
       MDDR_RAS_N,
       MDDR_ODT,
       MDDR_DQS_TMATCH_0_OUT,
       MDDR_DQS_TMATCH_0_IN,
       MDDR_CS_N,
       MDDR_CKE,
       MDDR_CAS_N,
       I2C_1_SDA,
       I2C_1_SCL,
       I2C_0_SDA,
       I2C_0_SCL,
       GPIO_3_M2F_c,
       GPIO_2_M2F_c,
       M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F,
       GPIO_1_M2F_c,
       GPIO_0_M2F_c,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE,
       CORECONFIGP_0_MDDR_APBmslave_PREADY,
       CORECONFIGP_0_MDDR_APBmslave_PSLVERR,
       CORECONFIGP_0_SOFT_M3_RESET_i_0,
       FAB_CCC_LOCK_c,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR,
       CORECONFIGP_0_SOFT_RESET_F2M_i_0,
       FAB_CCC_GL0_c,
       CORECONFIGP_0_MDDR_APBmslave_PENABLE,
       CORECONFIGP_0_MDDR_APBmslave_PSELx,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE,
       MDDR_CLK_N,
       MDDR_CLK
    );
inout  [7:0] MDDR_DQ;
inout  [0:0] MDDR_DM_RDQS;
output [2:0] MDDR_BA;
output [15:0] MDDR_ADDR;
output [15:2] M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR;
output [31:0] M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA;
output [15:0] CORECONFIGP_0_MDDR_APBmslave_PRDATA;
input  [31:0] M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA;
input  [10:2] M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR;
input  [15:0] M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA;
inout  [0:0] MDDR_DQS_N;
inout  [0:0] MDDR_DQS;
output FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA;
output MSS_ADLIB_INST_RNI7K43;
output un1_M2S_MSS_sb_0_4_i_0;
inout  SPI_1_SS0;
output SPI_1_DO;
input  SPI_1_DI;
inout  SPI_1_CLK;
inout  SPI_0_SS0;
output SPI_0_DO;
input  SPI_0_DI;
inout  SPI_0_CLK;
output MMUART_1_TXD;
input  MMUART_1_RXD;
output MMUART_0_TXD;
input  MMUART_0_RXD;
output MDDR_WE_N;
output MDDR_RESET_N;
output MDDR_RAS_N;
output MDDR_ODT;
output MDDR_DQS_TMATCH_0_OUT;
input  MDDR_DQS_TMATCH_0_IN;
output MDDR_CS_N;
output MDDR_CKE;
output MDDR_CAS_N;
inout  I2C_1_SDA;
inout  I2C_1_SCL;
inout  I2C_0_SDA;
inout  I2C_0_SCL;
output GPIO_3_M2F_c;
output GPIO_2_M2F_c;
output M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F;
output GPIO_1_M2F_c;
output GPIO_0_M2F_c;
output M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE;
output M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx;
output M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE;
output CORECONFIGP_0_MDDR_APBmslave_PREADY;
output CORECONFIGP_0_MDDR_APBmslave_PSLVERR;
input  CORECONFIGP_0_SOFT_M3_RESET_i_0;
input  FAB_CCC_LOCK_c;
input  M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY;
input  M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR;
input  CORECONFIGP_0_SOFT_RESET_F2M_i_0;
input  FAB_CCC_GL0_c;
input  CORECONFIGP_0_MDDR_APBmslave_PENABLE;
input  CORECONFIGP_0_MDDR_APBmslave_PSELx;
input  M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE;
output MDDR_CLK_N;
output MDDR_CLK;

    wire FIC_2_APB_M_PCLK, CONFIG_PRESET_N, SPI_1_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT, 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE, 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT, 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE, SPI_1_DI_PAD_Y, 
        SPI_1_CLK_PAD_Y, MSS_ADLIB_INST_SPI1_SCK_OUT, 
        MSS_ADLIB_INST_SPI1_SCK_OE, SPI_0_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, SPI_0_DI_PAD_Y, 
        SPI_0_CLK_PAD_Y, MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, 
        MMUART_0_RXD_PAD_Y, MSS_ADLIB_INST_DRAM_WEN, 
        MSS_ADLIB_INST_DRAM_RSTN, MSS_ADLIB_INST_DRAM_RASN, 
        MSS_ADLIB_INST_DRAM_ODT, \DRAM_FIFO_WE_OUT_net_0[0] , 
        MDDR_DQS_TMATCH_0_IN_PAD_Y, MDDR_DQ_7_PAD_Y, 
        \DRAM_DQ_OUT_net_0[7] , \DRAM_DQ_OE_net_0[7] , MDDR_DQ_6_PAD_Y, 
        \DRAM_DQ_OUT_net_0[6] , \DRAM_DQ_OE_net_0[6] , MDDR_DQ_5_PAD_Y, 
        \DRAM_DQ_OUT_net_0[5] , \DRAM_DQ_OE_net_0[5] , MDDR_DQ_4_PAD_Y, 
        \DRAM_DQ_OUT_net_0[4] , \DRAM_DQ_OE_net_0[4] , MDDR_DQ_3_PAD_Y, 
        \DRAM_DQ_OUT_net_0[3] , \DRAM_DQ_OE_net_0[3] , MDDR_DQ_2_PAD_Y, 
        \DRAM_DQ_OUT_net_0[2] , \DRAM_DQ_OE_net_0[2] , MDDR_DQ_1_PAD_Y, 
        \DRAM_DQ_OUT_net_0[1] , \DRAM_DQ_OE_net_0[1] , MDDR_DQ_0_PAD_Y, 
        \DRAM_DQ_OUT_net_0[0] , \DRAM_DQ_OE_net_0[0] , 
        MDDR_DM_RDQS_0_PAD_Y, \DRAM_DM_RDQS_OUT_net_0[0] , 
        \DM_OE_net_0[0] , MSS_ADLIB_INST_DRAM_CSN, 
        MSS_ADLIB_INST_DRAM_CKE, MSS_ADLIB_INST_DRAM_CASN, 
        \DRAM_BA_net_0[2] , \DRAM_BA_net_0[1] , \DRAM_BA_net_0[0] , 
        \DRAM_ADDR_net_0[15] , \DRAM_ADDR_net_0[14] , 
        \DRAM_ADDR_net_0[13] , \DRAM_ADDR_net_0[12] , 
        \DRAM_ADDR_net_0[11] , \DRAM_ADDR_net_0[10] , 
        \DRAM_ADDR_net_0[9] , \DRAM_ADDR_net_0[8] , 
        \DRAM_ADDR_net_0[7] , \DRAM_ADDR_net_0[6] , 
        \DRAM_ADDR_net_0[5] , \DRAM_ADDR_net_0[4] , 
        \DRAM_ADDR_net_0[3] , \DRAM_ADDR_net_0[2] , 
        \DRAM_ADDR_net_0[1] , \DRAM_ADDR_net_0[0] , I2C_1_SDA_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, I2C_1_SCL_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, I2C_0_SDA_PAD_Y, 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT, 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE, 
        I2C_0_SCL_PAD_Y, 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT, 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE, VCC_net_1, 
        GND_net_1, MDDR_DQS_0_PAD_Y, MSS_ADLIB_INST_DRAM_CLK, 
        \DRAM_DQS_OUT_net_0[0] , \DRAM_DQS_OE_net_0[0] ;
    
    INBUF #( .IOSTD("") )  MMUART_0_RXD_PAD (.PAD(MMUART_0_RXD), .Y(
        MMUART_0_RXD_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_6_PAD (.D(
        \DRAM_ADDR_net_0[6] ), .PAD(MDDR_ADDR[6]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_CAS_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_CASN), .PAD(MDDR_CAS_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_RESET_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_RSTN), .PAD(MDDR_RESET_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ODT_PAD (.D(
        MSS_ADLIB_INST_DRAM_ODT), .PAD(MDDR_ODT));
    CLKINT MSS_ADLIB_INST_RNI7K43_inst_1 (.A(CONFIG_PRESET_N), .Y(
        MSS_ADLIB_INST_RNI7K43));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_11_PAD (.D(
        \DRAM_ADDR_net_0[11] ), .PAD(MDDR_ADDR[11]));
    TRIBUFF MMUART_1_TXD_PAD (.D(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT), .E(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE), .PAD(
        MMUART_1_TXD));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_1_PAD (.PAD(MDDR_DQ[1]), .D(
        \DRAM_DQ_OUT_net_0[1] ), .E(\DRAM_DQ_OE_net_0[1] ), .Y(
        MDDR_DQ_1_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_7_PAD (.D(
        \DRAM_ADDR_net_0[7] ), .PAD(MDDR_ADDR[7]));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_3_PAD (.PAD(MDDR_DQ[3]), .D(
        \DRAM_DQ_OUT_net_0[3] ), .E(\DRAM_DQ_OE_net_0[3] ), .Y(
        MDDR_DQ_3_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_0_PAD (.PAD(MDDR_DQ[0]), .D(
        \DRAM_DQ_OUT_net_0[0] ), .E(\DRAM_DQ_OE_net_0[0] ), .Y(
        MDDR_DQ_0_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_12_PAD (.D(
        \DRAM_ADDR_net_0[12] ), .PAD(MDDR_ADDR[12]));
    VCC VCC (.Y(VCC_net_1));
    BIBUF SPI_1_SS0_PAD (.PAD(SPI_1_SS0), .D(
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT), .E(
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE), .Y(SPI_1_SS0_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_2_PAD (.PAD(MDDR_DQ[2]), .D(
        \DRAM_DQ_OUT_net_0[2] ), .E(\DRAM_DQ_OE_net_0[2] ), .Y(
        MDDR_DQ_2_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_CKE_PAD (.D(
        MSS_ADLIB_INST_DRAM_CKE), .PAD(MDDR_CKE));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_2_PAD (.D(
        \DRAM_ADDR_net_0[2] ), .PAD(MDDR_ADDR[2]));
    CLKINT FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA_inst_1 (.A(
        FIC_2_APB_M_PCLK), .Y(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA));
    TRIBUFF MMUART_0_TXD_PAD (.D(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT), .E(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE), .PAD(
        MMUART_0_TXD));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_13_PAD (.D(
        \DRAM_ADDR_net_0[13] ), .PAD(MDDR_ADDR[13]));
    BIBUF I2C_1_SDA_PAD (.PAD(I2C_1_SDA), .D(
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT), .E(
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE), .Y(
        I2C_1_SDA_PAD_Y));
    BIBUF I2C_1_SCL_PAD (.PAD(I2C_1_SCL), .D(
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT), .E(
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE), .Y(
        I2C_1_SCL_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_5_PAD (.D(
        \DRAM_ADDR_net_0[5] ), .PAD(MDDR_ADDR[5]));
    TRIBUFF SPI_1_DO_PAD (.D(MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT), .E(
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE), .PAD(SPI_1_DO));
    TRIBUFF SPI_0_DO_PAD (.D(
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT), .E(
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE), .PAD(SPI_0_DO));
    BIBUF_DIFF #( .IOSTD("SSTL18I") )  MDDR_DQS_0_PAD (.D(
        \DRAM_DQS_OUT_net_0[0] ), .E(\DRAM_DQS_OE_net_0[0] ), .PADP(
        MDDR_DQS[0]), .PADN(MDDR_DQS_N[0]), .Y(MDDR_DQS_0_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DM_RDQS_0_PAD (.PAD(
        MDDR_DM_RDQS[0]), .D(\DRAM_DM_RDQS_OUT_net_0[0] ), .E(
        \DM_OE_net_0[0] ), .Y(MDDR_DM_RDQS_0_PAD_Y));
    INBUF #( .IOSTD("") )  SPI_1_DI_PAD (.PAD(SPI_1_DI), .Y(
        SPI_1_DI_PAD_Y));
    BIBUF I2C_0_SCL_PAD (.PAD(I2C_0_SCL), .D(
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT), .E(
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE), .Y(
        I2C_0_SCL_PAD_Y));
    GND GND (.Y(GND_net_1));
    INBUF #( .IOSTD("") )  SPI_0_DI_PAD (.PAD(SPI_0_DI), .Y(
        SPI_0_DI_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_9_PAD (.D(
        \DRAM_ADDR_net_0[9] ), .PAD(MDDR_ADDR[9]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_BA_2_PAD (.D(
        \DRAM_BA_net_0[2] ), .PAD(MDDR_BA[2]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_14_PAD (.D(
        \DRAM_ADDR_net_0[14] ), .PAD(MDDR_ADDR[14]));
    MSS_075 #( .INIT(1438'h00000401003612000000000000000036100080000000000000000000000000000000000012036100000000000000000001203610000000001004000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33F00020200E0864A560003FFFFE4000000000000400000000F0F01C00000002D814010842108421000001FE34001FF8000000400000000000EF1007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(332.0)
         )  MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(GPIO_3_M2F_c), 
        .CAN_TX_EBL_MGPIO4A_H2F_A(), .CAN_TX_EBL_MGPIO4A_H2F_B(), 
        .CAN_TXBUS_MGPIO2A_H2F_A(), .CAN_TXBUS_MGPIO2A_H2F_B(
        GPIO_2_M2F_c), .CLK_CONFIG_APB(FIC_2_APB_M_PCLK), .COMMS_INT(), 
        .CONFIG_PRESET_N(CONFIG_PRESET_N), .EDAC_ERROR({nc0, nc1, nc2, 
        nc3, nc4, nc5, nc6, nc7}), .F_FM0_RDATA({nc8, nc9, nc10, nc11, 
        nc12, nc13, nc14, nc15, nc16, nc17, nc18, nc19, nc20, nc21, 
        nc22, nc23, nc24, nc25, nc26, nc27, nc28, nc29, nc30, nc31, 
        nc32, nc33, nc34, nc35, nc36, nc37, nc38, nc39}), 
        .F_FM0_READYOUT(), .F_FM0_RESP(), .F_HM0_ADDR({nc40, nc41, 
        nc42, nc43, nc44, nc45, nc46, nc47, nc48, nc49, nc50, nc51, 
        nc52, nc53, nc54, nc55, nc56, nc57, nc58, nc59, nc60, nc61, 
        nc62, nc63, nc64, nc65, nc66, nc67, nc68, nc69, nc70, nc71}), 
        .F_HM0_ENABLE(), .F_HM0_SEL(), .F_HM0_SIZE({nc72, nc73}), 
        .F_HM0_TRANS1(), .F_HM0_WDATA({nc74, nc75, nc76, nc77, nc78, 
        nc79, nc80, nc81, nc82, nc83, nc84, nc85, nc86, nc87, nc88, 
        nc89, nc90, nc91, nc92, nc93, nc94, nc95, nc96, nc97, nc98, 
        nc99, nc100, nc101, nc102, nc103, nc104, nc105}), .F_HM0_WRITE(
        ), .FAB_CHRGVBUS(), .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), 
        .FAB_DPPULLDOWN(), .FAB_DRVVBUS(), .FAB_IDPULLUP(), 
        .FAB_OPMODE({nc106, nc107}), .FAB_SUSPENDM(), .FAB_TERMSEL(), 
        .FAB_TXVALID(), .FAB_VCONTROL({nc108, nc109, nc110, nc111}), 
        .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({nc112, nc113}), 
        .FAB_XDATAOUT({nc114, nc115, nc116, nc117, nc118, nc119, nc120, 
        nc121}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc122, nc123}), 
        .FIC32_1_MASTER({nc124, nc125}), .FPGA_RESET_N(
        M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F), .GTX_CLK(), 
        .H2F_INTERRUPT({nc126, nc127, nc128, nc129, nc130, nc131, 
        nc132, nc133, nc134, nc135, nc136, nc137, nc138, nc139, nc140, 
        nc141}), .H2F_NMI(), .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(GPIO_1_M2F_c), .I2C1_SDA_MGPIO0A_H2F_A(
        ), .I2C1_SDA_MGPIO0A_H2F_B(GPIO_0_M2F_c), .MDCF(), .MDOENF(), 
        .MDOF(), .MMUART0_CTS_MGPIO19B_H2F_A(), 
        .MMUART0_CTS_MGPIO19B_H2F_B(), .MMUART0_DCD_MGPIO22B_H2F_A(), 
        .MMUART0_DCD_MGPIO22B_H2F_B(), .MMUART0_DSR_MGPIO20B_H2F_A(), 
        .MMUART0_DSR_MGPIO20B_H2F_B(), .MMUART0_DTR_MGPIO18B_H2F_A(), 
        .MMUART0_DTR_MGPIO18B_H2F_B(), .MMUART0_RI_MGPIO21B_H2F_A(), 
        .MMUART0_RI_MGPIO21B_H2F_B(), .MMUART0_RTS_MGPIO17B_H2F_A(), 
        .MMUART0_RTS_MGPIO17B_H2F_B(), .MMUART0_RXD_MGPIO28B_H2F_A(), 
        .MMUART0_RXD_MGPIO28B_H2F_B(), .MMUART0_SCK_MGPIO29B_H2F_A(), 
        .MMUART0_SCK_MGPIO29B_H2F_B(), .MMUART0_TXD_MGPIO27B_H2F_A(), 
        .MMUART0_TXD_MGPIO27B_H2F_B(), .MMUART1_DTR_MGPIO12B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_B(), 
        .MMUART1_RXD_MGPIO26B_H2F_A(), .MMUART1_RXD_MGPIO26B_H2F_B(), 
        .MMUART1_SCK_MGPIO25B_H2F_A(), .MMUART1_SCK_MGPIO25B_H2F_B(), 
        .MMUART1_TXD_MGPIO24B_H2F_A(), .MMUART1_TXD_MGPIO24B_H2F_B(), 
        .MPLL_LOCK(), .PER2_FABRIC_PADDR({
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[14], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[11], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]}), 
        .PER2_FABRIC_PENABLE(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE), 
        .PER2_FABRIC_PSEL(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx), 
        .PER2_FABRIC_PWDATA({
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[31], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[30], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[29], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[28], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[27], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[26], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[25], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[24], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[23], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[22], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[21], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[20], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[19], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[18], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[17], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]}), 
        .PER2_FABRIC_PWRITE(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE), .RTC_MATCH(), 
        .SLEEPDEEP(), .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), 
        .SMBALERT_NO1(), .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc142, nc143, nc144, nc145, 
        nc146, nc147, nc148, nc149, nc150, nc151}), .TRACECLK(), 
        .TRACEDATA({nc152, nc153, nc154, nc155}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc156, nc157, nc158, 
        nc159}), .TXDF({nc160, nc161, nc162, nc163, nc164, nc165, 
        nc166, nc167}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc168, nc169, nc170, nc171})
        , .F_BRESP_HRESP0({nc172, nc173}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc174, nc175, nc176, nc177, nc178, nc179, 
        nc180, nc181, nc182, nc183, nc184, nc185, nc186, nc187, nc188, 
        nc189, nc190, nc191, nc192, nc193, nc194, nc195, nc196, nc197, 
        nc198, nc199, nc200, nc201, nc202, nc203, nc204, nc205, nc206, 
        nc207, nc208, nc209, nc210, nc211, nc212, nc213, nc214, nc215, 
        nc216, nc217, nc218, nc219, nc220, nc221, nc222, nc223, nc224, 
        nc225, nc226, nc227, nc228, nc229, nc230, nc231, nc232, nc233, 
        nc234, nc235, nc236, nc237}), .F_RID({nc238, nc239, nc240, 
        nc241}), .F_RLAST(), .F_RRESP_HRESP1({nc242, nc243}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[15], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[14], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[13], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[12], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[11], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[10], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[9], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[8], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[7], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[6], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[5], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[4], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[3], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[2], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[1], 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]}), .MDDR_FABRIC_PREADY(
        CORECONFIGP_0_MDDR_APBmslave_PREADY), .MDDR_FABRIC_PSLVERR(
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR), .CAN_RXBUS_F2H_SCP(
        VCC_net_1), .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(
        VCC_net_1), .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({
        VCC_net_1, VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), .F2HCALIB(
        VCC_net_1), .F_DMAREADY({VCC_net_1, VCC_net_1}), .F_FM0_ADDR({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_FM0_ENABLE(GND_net_1), 
        .F_FM0_MASTLOCK(GND_net_1), .F_FM0_READY(VCC_net_1), 
        .F_FM0_SEL(GND_net_1), .F_FM0_SIZE({GND_net_1, GND_net_1}), 
        .F_FM0_TRANS1(GND_net_1), .F_FM0_WDATA({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_FM0_WRITE(GND_net_1), .F_HM0_RDATA({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_HM0_READY(VCC_net_1), .F_HM0_RESP(GND_net_1), .FAB_AVALID(
        VCC_net_1), .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(VCC_net_1), 
        .FAB_LINESTATE({VCC_net_1, VCC_net_1}), .FAB_M3_RESET_N(
        CORECONFIGP_0_SOFT_M3_RESET_i_0), .FAB_PLL_LOCK(FAB_CCC_LOCK_c)
        , .FAB_RXACTIVE(VCC_net_1), .FAB_RXERROR(VCC_net_1), 
        .FAB_RXVALID(VCC_net_1), .FAB_RXVALIDH(GND_net_1), 
        .FAB_SESSEND(VCC_net_1), .FAB_TXREADY(VCC_net_1), 
        .FAB_VBUSVALID(VCC_net_1), .FAB_VSTATUS({VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .FAB_XDATAIN({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .GTX_CLKPF(VCC_net_1), .I2C0_BCLK(VCC_net_1), 
        .I2C0_SCL_F2H_SCP(VCC_net_1), .I2C0_SDA_F2H_SCP(VCC_net_1), 
        .I2C1_BCLK(VCC_net_1), .I2C1_SCL_F2H_SCP(VCC_net_1), 
        .I2C1_SDA_F2H_SCP(VCC_net_1), .MDIF(VCC_net_1), 
        .MGPIO0A_F2H_GPIN(VCC_net_1), .MGPIO10A_F2H_GPIN(VCC_net_1), 
        .MGPIO11A_F2H_GPIN(VCC_net_1), .MGPIO11B_F2H_GPIN(VCC_net_1), 
        .MGPIO12A_F2H_GPIN(VCC_net_1), .MGPIO13A_F2H_GPIN(VCC_net_1), 
        .MGPIO14A_F2H_GPIN(VCC_net_1), .MGPIO15A_F2H_GPIN(VCC_net_1), 
        .MGPIO16A_F2H_GPIN(VCC_net_1), .MGPIO17B_F2H_GPIN(VCC_net_1), 
        .MGPIO18B_F2H_GPIN(VCC_net_1), .MGPIO19B_F2H_GPIN(VCC_net_1), 
        .MGPIO1A_F2H_GPIN(VCC_net_1), .MGPIO20B_F2H_GPIN(VCC_net_1), 
        .MGPIO21B_F2H_GPIN(VCC_net_1), .MGPIO22B_F2H_GPIN(VCC_net_1), 
        .MGPIO24B_F2H_GPIN(VCC_net_1), .MGPIO25B_F2H_GPIN(VCC_net_1), 
        .MGPIO26B_F2H_GPIN(VCC_net_1), .MGPIO27B_F2H_GPIN(VCC_net_1), 
        .MGPIO28B_F2H_GPIN(VCC_net_1), .MGPIO29B_F2H_GPIN(VCC_net_1), 
        .MGPIO2A_F2H_GPIN(VCC_net_1), .MGPIO30B_F2H_GPIN(VCC_net_1), 
        .MGPIO31B_F2H_GPIN(VCC_net_1), .MGPIO3A_F2H_GPIN(VCC_net_1), 
        .MGPIO4A_F2H_GPIN(VCC_net_1), .MGPIO5A_F2H_GPIN(VCC_net_1), 
        .MGPIO6A_F2H_GPIN(VCC_net_1), .MGPIO7A_F2H_GPIN(VCC_net_1), 
        .MGPIO8A_F2H_GPIN(VCC_net_1), .MGPIO9A_F2H_GPIN(VCC_net_1), 
        .MMUART0_CTS_F2H_SCP(VCC_net_1), .MMUART0_DCD_F2H_SCP(
        VCC_net_1), .MMUART0_DSR_F2H_SCP(VCC_net_1), 
        .MMUART0_DTR_F2H_SCP(VCC_net_1), .MMUART0_RI_F2H_SCP(VCC_net_1)
        , .MMUART0_RTS_F2H_SCP(VCC_net_1), .MMUART0_RXD_F2H_SCP(
        VCC_net_1), .MMUART0_SCK_F2H_SCP(VCC_net_1), 
        .MMUART0_TXD_F2H_SCP(VCC_net_1), .MMUART1_CTS_F2H_SCP(
        VCC_net_1), .MMUART1_DCD_F2H_SCP(VCC_net_1), 
        .MMUART1_DSR_F2H_SCP(VCC_net_1), .MMUART1_RI_F2H_SCP(VCC_net_1)
        , .MMUART1_RTS_F2H_SCP(VCC_net_1), .MMUART1_RXD_F2H_SCP(
        VCC_net_1), .MMUART1_SCK_F2H_SCP(VCC_net_1), 
        .MMUART1_TXD_F2H_SCP(VCC_net_1), .PER2_FABRIC_PRDATA({
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[31], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[30], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[29], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[28], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[27], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[26], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[25], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[24], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[23], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[22], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[21], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[20], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[19], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[18], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1], 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]}), 
        .PER2_FABRIC_PREADY(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY), 
        .PER2_FABRIC_PSLVERR(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR), .RCGF({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .RX_CLKPF(VCC_net_1), .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), 
        .RX_EV(VCC_net_1), .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .SLEEPHOLDREQ(GND_net_1), .SMBALERT_NI0(VCC_net_1), 
        .SMBALERT_NI1(VCC_net_1), .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(
        VCC_net_1), .SPI0_CLK_IN(VCC_net_1), .SPI0_SDI_F2H_SCP(
        VCC_net_1), .SPI0_SDO_F2H_SCP(VCC_net_1), .SPI0_SS0_F2H_SCP(
        VCC_net_1), .SPI0_SS1_F2H_SCP(VCC_net_1), .SPI0_SS2_F2H_SCP(
        VCC_net_1), .SPI0_SS3_F2H_SCP(VCC_net_1), .SPI1_CLK_IN(
        VCC_net_1), .SPI1_SDI_F2H_SCP(VCC_net_1), .SPI1_SDO_F2H_SCP(
        VCC_net_1), .SPI1_SS0_F2H_SCP(VCC_net_1), .SPI1_SS1_F2H_SCP(
        VCC_net_1), .SPI1_SS2_F2H_SCP(VCC_net_1), .SPI1_SS3_F2H_SCP(
        VCC_net_1), .TX_CLKPF(VCC_net_1), .USER_MSS_GPIO_RESET_N(
        VCC_net_1), .USER_MSS_RESET_N(CORECONFIGP_0_SOFT_RESET_F2M_i_0)
        , .XCLK_FAB(VCC_net_1), .CLK_BASE(FAB_CCC_GL0_c), 
        .CLK_MDDR_APB(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), 
        .F_ARADDR_HADDR1({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .F_ARBURST_HTRANS1({
        GND_net_1, GND_net_1}), .F_ARID_HSEL1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLEN_HBURST1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLOCK_HMASTLOCK1({GND_net_1, 
        GND_net_1}), .F_ARSIZE_HSIZE1({GND_net_1, GND_net_1}), 
        .F_ARVALID_HWRITE1(GND_net_1), .F_AWADDR_HADDR0({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_AWBURST_HTRANS0({GND_net_1, GND_net_1}), 
        .F_AWID_HSEL0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLEN_HBURST0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLOCK_HMASTLOCK0({GND_net_1, GND_net_1}), .F_AWSIZE_HSIZE0({
        GND_net_1, GND_net_1}), .F_AWVALID_HWRITE0(GND_net_1), 
        .F_BREADY(GND_net_1), .F_RMW_AXI(GND_net_1), .F_RREADY(
        GND_net_1), .F_WDATA_HWDATA01({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_WID_HREADY01({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_WLAST(GND_net_1), .F_WSTRB({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_WVALID(GND_net_1), 
        .FPGA_MDDR_ARESET_N(VCC_net_1), .MDDR_FABRIC_PADDR({
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[2]}), .MDDR_FABRIC_PENABLE(
        CORECONFIGP_0_MDDR_APBmslave_PENABLE), .MDDR_FABRIC_PSEL(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .MDDR_FABRIC_PWDATA({
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[15], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[14], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[13], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[12], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[11], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[2], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[1], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[0]}), .MDDR_FABRIC_PWRITE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE), .PRESET_N(
        MSS_ADLIB_INST_RNI7K43), .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(
        GND_net_1), .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, MDDR_DM_RDQS_0_PAD_Y}), .DRAM_DQ_IN({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, MDDR_DQ_7_PAD_Y, 
        MDDR_DQ_6_PAD_Y, MDDR_DQ_5_PAD_Y, MDDR_DQ_4_PAD_Y, 
        MDDR_DQ_3_PAD_Y, MDDR_DQ_2_PAD_Y, MDDR_DQ_1_PAD_Y, 
        MDDR_DQ_0_PAD_Y}), .DRAM_DQS_IN({GND_net_1, GND_net_1, 
        MDDR_DQS_0_PAD_Y}), .DRAM_FIFO_WE_IN({GND_net_1, 
        MDDR_DQS_TMATCH_0_IN_PAD_Y}), .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(
        I2C_0_SCL_PAD_Y), .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(
        I2C_0_SDA_PAD_Y), .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(
        I2C_1_SCL_PAD_Y), .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(
        I2C_1_SDA_PAD_Y), .MGPIO0B_IN(GND_net_1), .MGPIO10B_IN(
        GND_net_1), .MGPIO1B_IN(GND_net_1), .MGPIO25A_IN(GND_net_1), 
        .MGPIO26A_IN(GND_net_1), .MGPIO27A_IN(GND_net_1), .MGPIO28A_IN(
        GND_net_1), .MGPIO29A_IN(GND_net_1), .MGPIO2B_IN(GND_net_1), 
        .MGPIO30A_IN(GND_net_1), .MGPIO31A_IN(GND_net_1), .MGPIO3B_IN(
        GND_net_1), .MGPIO4B_IN(GND_net_1), .MGPIO5B_IN(GND_net_1), 
        .MGPIO6B_IN(GND_net_1), .MGPIO7B_IN(GND_net_1), .MGPIO8B_IN(
        GND_net_1), .MGPIO9B_IN(GND_net_1), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND_net_1), 
        .MMUART0_DCD_MGPIO22B_IN(GND_net_1), .MMUART0_DSR_MGPIO20B_IN(
        GND_net_1), .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND_net_1), 
        .MMUART0_RI_MGPIO21B_IN(GND_net_1), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(MMUART_0_RXD_PAD_Y), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_CTS_MGPIO13B_IN(GND_net_1), .MMUART1_DCD_MGPIO16B_IN(
        GND_net_1), .MMUART1_DSR_MGPIO14B_IN(GND_net_1), 
        .MMUART1_DTR_MGPIO12B_IN(GND_net_1), .MMUART1_RI_MGPIO15B_IN(
        GND_net_1), .MMUART1_RTS_MGPIO11B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(MMUART_1_RXD_PAD_Y), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        SPI_0_CLK_PAD_Y), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(SPI_0_DI_PAD_Y)
        , .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(SPI_0_SS0_PAD_Y), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND_net_1), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND_net_1), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND_net_1), 
        .SPI0_SS4_MGPIO19A_IN(GND_net_1), .SPI0_SS5_MGPIO20A_IN(
        GND_net_1), .SPI0_SS6_MGPIO21A_IN(GND_net_1), 
        .SPI0_SS7_MGPIO22A_IN(GND_net_1), .SPI1_SCK_IN(SPI_1_CLK_PAD_Y)
        , .SPI1_SDI_MGPIO11A_IN(SPI_1_DI_PAD_Y), .SPI1_SDO_MGPIO12A_IN(
        GND_net_1), .SPI1_SS0_MGPIO13A_IN(SPI_1_SS0_PAD_Y), 
        .SPI1_SS1_MGPIO14A_IN(GND_net_1), .SPI1_SS2_MGPIO15A_IN(
        GND_net_1), .SPI1_SS3_MGPIO16A_IN(GND_net_1), 
        .SPI1_SS4_MGPIO17A_IN(GND_net_1), .SPI1_SS5_MGPIO18A_IN(
        GND_net_1), .SPI1_SS6_MGPIO23A_IN(GND_net_1), 
        .SPI1_SS7_MGPIO24A_IN(GND_net_1), .USBC_XCLK_IN(GND_net_1), 
        .USBD_DATA0_IN(GND_net_1), .USBD_DATA1_IN(GND_net_1), 
        .USBD_DATA2_IN(GND_net_1), .USBD_DATA3_IN(GND_net_1), 
        .USBD_DATA4_IN(GND_net_1), .USBD_DATA5_IN(GND_net_1), 
        .USBD_DATA6_IN(GND_net_1), .USBD_DATA7_MGPIO23B_IN(GND_net_1), 
        .USBD_DIR_IN(GND_net_1), .USBD_NXT_IN(GND_net_1), .USBD_STP_IN(
        GND_net_1), .USBD_XCLK_IN(GND_net_1), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({
        \DRAM_ADDR_net_0[15] , \DRAM_ADDR_net_0[14] , 
        \DRAM_ADDR_net_0[13] , \DRAM_ADDR_net_0[12] , 
        \DRAM_ADDR_net_0[11] , \DRAM_ADDR_net_0[10] , 
        \DRAM_ADDR_net_0[9] , \DRAM_ADDR_net_0[8] , 
        \DRAM_ADDR_net_0[7] , \DRAM_ADDR_net_0[6] , 
        \DRAM_ADDR_net_0[5] , \DRAM_ADDR_net_0[4] , 
        \DRAM_ADDR_net_0[3] , \DRAM_ADDR_net_0[2] , 
        \DRAM_ADDR_net_0[1] , \DRAM_ADDR_net_0[0] }), .DRAM_BA({
        \DRAM_BA_net_0[2] , \DRAM_BA_net_0[1] , \DRAM_BA_net_0[0] }), 
        .DRAM_CASN(MSS_ADLIB_INST_DRAM_CASN), .DRAM_CKE(
        MSS_ADLIB_INST_DRAM_CKE), .DRAM_CLK(MSS_ADLIB_INST_DRAM_CLK), 
        .DRAM_CSN(MSS_ADLIB_INST_DRAM_CSN), .DRAM_DM_RDQS_OUT({nc244, 
        nc245, \DRAM_DM_RDQS_OUT_net_0[0] }), .DRAM_DQ_OUT({nc246, 
        nc247, nc248, nc249, nc250, nc251, nc252, nc253, nc254, nc255, 
        \DRAM_DQ_OUT_net_0[7] , \DRAM_DQ_OUT_net_0[6] , 
        \DRAM_DQ_OUT_net_0[5] , \DRAM_DQ_OUT_net_0[4] , 
        \DRAM_DQ_OUT_net_0[3] , \DRAM_DQ_OUT_net_0[2] , 
        \DRAM_DQ_OUT_net_0[1] , \DRAM_DQ_OUT_net_0[0] }), 
        .DRAM_DQS_OUT({nc256, nc257, \DRAM_DQS_OUT_net_0[0] }), 
        .DRAM_FIFO_WE_OUT({nc258, \DRAM_FIFO_WE_OUT_net_0[0] }), 
        .DRAM_ODT(MSS_ADLIB_INST_DRAM_ODT), .DRAM_RASN(
        MSS_ADLIB_INST_DRAM_RASN), .DRAM_RSTN(MSS_ADLIB_INST_DRAM_RSTN)
        , .DRAM_WEN(MSS_ADLIB_INST_DRAM_WEN), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT), .MGPIO0B_OUT()
        , .MGPIO10B_OUT(), .MGPIO1B_OUT(), .MGPIO25A_OUT(), 
        .MGPIO26A_OUT(), .MGPIO27A_OUT(), .MGPIO28A_OUT(), 
        .MGPIO29A_OUT(), .MGPIO2B_OUT(), .MGPIO30A_OUT(), 
        .MGPIO31A_OUT(), .MGPIO3B_OUT(), .MGPIO4B_OUT(), .MGPIO5B_OUT()
        , .MGPIO6B_OUT(), .MGPIO7B_OUT(), .MGPIO8B_OUT(), .MGPIO9B_OUT(
        ), .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT), 
        .MMUART1_CTS_MGPIO13B_OUT(), .MMUART1_DCD_MGPIO16B_OUT(), 
        .MMUART1_DSR_MGPIO14B_OUT(), .MMUART1_DTR_MGPIO12B_OUT(), 
        .MMUART1_RI_MGPIO15B_OUT(), .MMUART1_RTS_MGPIO11B_OUT(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI0_SS4_MGPIO19A_OUT(), 
        .SPI0_SS5_MGPIO20A_OUT(), .SPI0_SS6_MGPIO21A_OUT(), 
        .SPI0_SS7_MGPIO22A_OUT(), .SPI1_SCK_OUT(
        MSS_ADLIB_INST_SPI1_SCK_OUT), .SPI1_SDI_MGPIO11A_OUT(), 
        .SPI1_SDO_MGPIO12A_OUT(MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT), 
        .SPI1_SS0_MGPIO13A_OUT(MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT), 
        .SPI1_SS1_MGPIO14A_OUT(), .SPI1_SS2_MGPIO15A_OUT(), 
        .SPI1_SS3_MGPIO16A_OUT(), .SPI1_SS4_MGPIO17A_OUT(), 
        .SPI1_SS5_MGPIO18A_OUT(), .SPI1_SS6_MGPIO23A_OUT(), 
        .SPI1_SS7_MGPIO24A_OUT(), .USBC_XCLK_OUT(), .USBD_DATA0_OUT(), 
        .USBD_DATA1_OUT(), .USBD_DATA2_OUT(), .USBD_DATA3_OUT(), 
        .USBD_DATA4_OUT(), .USBD_DATA5_OUT(), .USBD_DATA6_OUT(), 
        .USBD_DATA7_MGPIO23B_OUT(), .USBD_DIR_OUT(), .USBD_NXT_OUT(), 
        .USBD_STP_OUT(), .USBD_XCLK_OUT(), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc259, nc260, 
        \DM_OE_net_0[0] }), .DRAM_DQ_OE({nc261, nc262, nc263, nc264, 
        nc265, nc266, nc267, nc268, nc269, nc270, 
        \DRAM_DQ_OE_net_0[7] , \DRAM_DQ_OE_net_0[6] , 
        \DRAM_DQ_OE_net_0[5] , \DRAM_DQ_OE_net_0[4] , 
        \DRAM_DQ_OE_net_0[3] , \DRAM_DQ_OE_net_0[2] , 
        \DRAM_DQ_OE_net_0[1] , \DRAM_DQ_OE_net_0[0] }), .DRAM_DQS_OE({
        nc271, nc272, \DRAM_DQS_OE_net_0[0] }), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE), .MGPIO0B_OE(), 
        .MGPIO10B_OE(), .MGPIO1B_OE(), .MGPIO25A_OE(), .MGPIO26A_OE(), 
        .MGPIO27A_OE(), .MGPIO28A_OE(), .MGPIO29A_OE(), .MGPIO2B_OE(), 
        .MGPIO30A_OE(), .MGPIO31A_OE(), .MGPIO3B_OE(), .MGPIO4B_OE(), 
        .MGPIO5B_OE(), .MGPIO6B_OE(), .MGPIO7B_OE(), .MGPIO8B_OE(), 
        .MGPIO9B_OE(), .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE), 
        .MMUART1_CTS_MGPIO13B_OE(), .MMUART1_DCD_MGPIO16B_OE(), 
        .MMUART1_DSR_MGPIO14B_OE(), .MMUART1_DTR_MGPIO12B_OE(), 
        .MMUART1_RI_MGPIO15B_OE(), .MMUART1_RTS_MGPIO11B_OE(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OE(
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI0_SS4_MGPIO19A_OE(), 
        .SPI0_SS5_MGPIO20A_OE(), .SPI0_SS6_MGPIO21A_OE(), 
        .SPI0_SS7_MGPIO22A_OE(), .SPI1_SCK_OE(
        MSS_ADLIB_INST_SPI1_SCK_OE), .SPI1_SDI_MGPIO11A_OE(), 
        .SPI1_SDO_MGPIO12A_OE(MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE), 
        .SPI1_SS0_MGPIO13A_OE(MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE), 
        .SPI1_SS1_MGPIO14A_OE(), .SPI1_SS2_MGPIO15A_OE(), 
        .SPI1_SS3_MGPIO16A_OE(), .SPI1_SS4_MGPIO17A_OE(), 
        .SPI1_SS5_MGPIO18A_OE(), .SPI1_SS6_MGPIO23A_OE(), 
        .SPI1_SS7_MGPIO24A_OE(), .USBC_XCLK_OE(), .USBD_DATA0_OE(), 
        .USBD_DATA1_OE(), .USBD_DATA2_OE(), .USBD_DATA3_OE(), 
        .USBD_DATA4_OE(), .USBD_DATA5_OE(), .USBD_DATA6_OE(), 
        .USBD_DATA7_MGPIO23B_OE(), .USBD_DIR_OE(), .USBD_NXT_OE(), 
        .USBD_STP_OE(), .USBD_XCLK_OE());
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_RAS_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_RASN), .PAD(MDDR_RAS_N));
    BIBUF SPI_0_CLK_PAD (.PAD(SPI_0_CLK), .D(
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT), .E(
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE), .Y(SPI_0_CLK_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_4_PAD (.PAD(MDDR_DQ[4]), .D(
        \DRAM_DQ_OUT_net_0[4] ), .E(\DRAM_DQ_OE_net_0[4] ), .Y(
        MDDR_DQ_4_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_10_PAD (.D(
        \DRAM_ADDR_net_0[10] ), .PAD(MDDR_ADDR[10]));
    BIBUF I2C_0_SDA_PAD (.PAD(I2C_0_SDA), .D(
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT), .E(
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE), .Y(
        I2C_0_SDA_PAD_Y));
    INBUF #( .IOSTD("SSTL18I") )  MDDR_DQS_TMATCH_0_IN_PAD (.PAD(
        MDDR_DQS_TMATCH_0_IN), .Y(MDDR_DQS_TMATCH_0_IN_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_CS_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_CSN), .PAD(MDDR_CS_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_4_PAD (.D(
        \DRAM_ADDR_net_0[4] ), .PAD(MDDR_ADDR[4]));
    BIBUF SPI_0_SS0_PAD (.PAD(SPI_0_SS0), .D(
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT), .E(
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE), .Y(
        SPI_0_SS0_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_7_PAD (.PAD(MDDR_DQ[7]), .D(
        \DRAM_DQ_OUT_net_0[7] ), .E(\DRAM_DQ_OE_net_0[7] ), .Y(
        MDDR_DQ_7_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_WE_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_WEN), .PAD(MDDR_WE_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_8_PAD (.D(
        \DRAM_ADDR_net_0[8] ), .PAD(MDDR_ADDR[8]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_15_PAD (.D(
        \DRAM_ADDR_net_0[15] ), .PAD(MDDR_ADDR[15]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_0_PAD (.D(
        \DRAM_ADDR_net_0[0] ), .PAD(MDDR_ADDR[0]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_1_PAD (.D(
        \DRAM_ADDR_net_0[1] ), .PAD(MDDR_ADDR[1]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_3_PAD (.D(
        \DRAM_ADDR_net_0[3] ), .PAD(MDDR_ADDR[3]));
    INBUF #( .IOSTD("") )  MMUART_1_RXD_PAD (.PAD(MMUART_1_RXD), .Y(
        MMUART_1_RXD_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_BA_0_PAD (.D(
        \DRAM_BA_net_0[0] ), .PAD(MDDR_BA[0]));
    CFG1 #( .INIT(2'h1) )  FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA_0 (
        .A(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .Y(
        un1_M2S_MSS_sb_0_4_i_0));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_6_PAD (.PAD(MDDR_DQ[6]), .D(
        \DRAM_DQ_OUT_net_0[6] ), .E(\DRAM_DQ_OE_net_0[6] ), .Y(
        MDDR_DQ_6_PAD_Y));
    OUTBUF_DIFF #( .IOSTD("SSTL18I") )  MDDR_CLK_PAD (.D(
        MSS_ADLIB_INST_DRAM_CLK), .PADP(MDDR_CLK), .PADN(MDDR_CLK_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_DQS_TMATCH_0_OUT_PAD (.D(
        \DRAM_FIFO_WE_OUT_net_0[0] ), .PAD(MDDR_DQS_TMATCH_0_OUT));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_BA_1_PAD (.D(
        \DRAM_BA_net_0[1] ), .PAD(MDDR_BA[1]));
    BIBUF SPI_1_CLK_PAD (.PAD(SPI_1_CLK), .D(
        MSS_ADLIB_INST_SPI1_SCK_OUT), .E(MSS_ADLIB_INST_SPI1_SCK_OE), 
        .Y(SPI_1_CLK_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_5_PAD (.PAD(MDDR_DQ[5]), .D(
        \DRAM_DQ_OUT_net_0[5] ), .E(\DRAM_DQ_OE_net_0[5] ), .Y(
        MDDR_DQ_5_PAD_Y));
    
endmodule


module M2S_MSS_sb_CCC_0_FCCC(
       FAB_CCC_GL0_c,
       FAB_CCC_LOCK_c,
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FAB_CCC_GL0_c;
output FAB_CCC_LOCK_c;
input  FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GL0_net, VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CLKINT GL0_INST (.A(GL0_net), .Y(FAB_CCC_GL0_c));
    CCC #( .INIT(210'h0000007FB8000044D74000318C6318C1F18C61EC0404040400301)
        , .VCOFREQUENCY(800.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(
        FAB_CCC_LOCK_c), .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), 
        .CLK2(VCC_net_1), .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), 
        .NGMUX1_SEL(GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(
        GND_net_1), .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(
        VCC_net_1), .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(
        VCC_net_1), .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(
        VCC_net_1), .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(
        VCC_net_1), .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(GL0_net), .GL1(), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), 
        .RCOSC_1MHZ(GND_net_1), .XTLOSC(GND_net_1));
    
endmodule


module CoreConfigP_Z1(
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA,
       CORECONFIGP_0_MDDR_APBmslave_PRDATA,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_6,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_7,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_8,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_9,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_10,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_12,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_0,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_1,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_2,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_3,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_4,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_5,
       CORECONFIGP_0_SOFT_RESET_F2M_i_0,
       CORECONFIGP_0_SOFT_M3_RESET_i_0,
       MSS_ADLIB_INST_RNI7K43,
       FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA,
       CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET,
       CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET,
       CORECONFIGP_0_CONFIG1_DONE,
       CORECONFIGP_0_CONFIG2_DONE,
       CORECONFIGP_0_SOFT_SDIF0_PHY_RESET,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE,
       un1_M2S_MSS_sb_0_4_i_0,
       INIT_DONE_int,
       CORERESETP_0_SDIF_RELEASED,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE,
       CORECONFIGP_0_MDDR_APBmslave_PENABLE,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx,
       M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE,
       CORECONFIGP_0_MDDR_APBmslave_PREADY,
       CORECONFIGP_0_MDDR_APBmslave_PSELx,
       N_39,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR,
       CORECONFIGP_0_MDDR_APBmslave_PSLVERR
    );
input  [15:2] M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR;
output [31:0] M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA;
input  [31:0] M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA;
output [31:0] M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA;
input  [31:0] M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA;
input  [15:0] CORECONFIGP_0_MDDR_APBmslave_PRDATA;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_6;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_7;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_8;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_9;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_10;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_12;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_0;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_1;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_2;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_3;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_4;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_5;
output CORECONFIGP_0_SOFT_RESET_F2M_i_0;
output CORECONFIGP_0_SOFT_M3_RESET_i_0;
input  MSS_ADLIB_INST_RNI7K43;
input  FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA;
output CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET;
output CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET;
output CORECONFIGP_0_CONFIG1_DONE;
output CORECONFIGP_0_CONFIG2_DONE;
output CORECONFIGP_0_SOFT_SDIF0_PHY_RESET;
output M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY;
output M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE;
input  M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE;
input  un1_M2S_MSS_sb_0_4_i_0;
input  INIT_DONE_int;
input  CORERESETP_0_SDIF_RELEASED;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE;
output CORECONFIGP_0_MDDR_APBmslave_PENABLE;
input  M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY;
input  M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx;
input  M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE;
input  CORECONFIGP_0_MDDR_APBmslave_PREADY;
output CORECONFIGP_0_MDDR_APBmslave_PSELx;
output N_39;
input  M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR;
input  CORECONFIGP_0_MDDR_APBmslave_PSLVERR;

    wire CORECONFIGP_0_SOFT_RESET_F2M, CORECONFIGP_0_SOFT_M3_RESET, 
        VCC_net_1, state_347_d, GND_net_1, 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] , 
        \soft_reset_reg[12]_net_1 , soft_reset_reg6, 
        \soft_reset_reg[13]_net_1 , \soft_reset_reg[14]_net_1 , 
        control_reg_15, \prdata[29] , \state[1]_net_1 , \prdata[30] , 
        \prdata[31] , \soft_reset_reg[0]_net_1 , 
        \soft_reset_reg[3]_net_1 , \soft_reset_reg[4]_net_1 , 
        \soft_reset_reg[5]_net_1 , \soft_reset_reg[6]_net_1 , 
        \soft_reset_reg[8]_net_1 , \soft_reset_reg[9]_net_1 , 
        \soft_reset_reg[10]_net_1 , \soft_reset_reg[11]_net_1 , 
        \prdata[14] , \prdata[15] , \prdata[16] , \prdata[17] , 
        \prdata[18] , \prdata[19] , \prdata[20] , \prdata[21] , 
        \prdata[22] , \prdata[23] , \prdata[24] , \prdata[25] , 
        \prdata[26] , \prdata[27] , \prdata[28] , \prdata[0] , 
        \prdata[1] , \prdata[2] , \prdata[3] , \prdata[4] , 
        \prdata[5] , \prdata[6] , \prdata[7] , \prdata[8] , 
        \prdata[9] , \prdata[10] , \prdata[11] , \prdata[12] , 
        \prdata[13] , N_51_i_0, pslverr, \state[0]_net_1 , 
        \state_ns[0] , \state_ns[1] , psel_net_1, state_347_d_i_0, 
        INIT_DONE_q1_net_1, SDIF_RELEASED_q1_net_1, INIT_DONE_q2_net_1, 
        SDIF_RELEASED_q2_net_1, N_16_i_0, MDDR_PENABLE_2, 
        prdata_0_iv_0_a3_out_0, prdata_0_iv_0_a2_1_out, g1_0_0_0, N_50, 
        N_46, \prdata_0_iv_0_a2_0[17] , soft_reset_reg6_0_a2_0_net_1, 
        control_reg_15_0_a2_0_net_1, N_48, \prdata_0_iv_0_a2_0[16] , 
        \prdata_0_iv_0_a2_1[5] , \prdata_0_iv_0_a2_1[0]_net_1 , N_38, 
        \prdata_0_iv_0_a2_1[1] , control_reg_15_4, N_113, N_126, N_122, 
        \prdata_0_iv_0_0[5]_net_1 , \prdata_0_iv_0_0[8]_net_1 , N_115, 
        \prdata_0_iv_0_0[1]_net_1 , \prdata_0_iv_0_0[14]_net_1 , 
        \prdata_0_iv_0_0[15]_net_1 , \prdata_0_iv_0_0[12]_net_1 , 
        \prdata_0_iv_0_0[13]_net_1 , \prdata_0_iv_0_0[10]_net_1 , 
        \prdata_0_iv_0_0[11]_net_1 , \prdata_0_iv_0_0[9]_net_1 , 
        \prdata_0_iv_0_0[6]_net_1 , \prdata_0_iv_0_0[7]_net_1 , 
        \prdata_0_iv_0_0[2]_net_1 , \prdata_0_iv_0_0[3]_net_1 , 
        \prdata_0_iv_0_0[4]_net_1 , \prdata_0_iv_0_tz[0]_net_1 , 
        \prdata_0_iv_0_0[0]_net_1 ;
    
    SLE \FIC_2_APB_M_PRDATA[13]  (.D(\prdata[13] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]));
    SLE \state[0]  (.D(\state_ns[0] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(VCC_net_1), .ALn(
        MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[0]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \prdata_0_iv_0_tz[0]  (.A(
        prdata_0_iv_0_a3_out_0), .B(\soft_reset_reg[0]_net_1 ), .C(
        \prdata_0_iv_0_a2_1[0]_net_1 ), .D(prdata_0_iv_0_a2_1_out), .Y(
        \prdata_0_iv_0_tz[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[27]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[27]), .Y(\prdata[27] ));
    SLE \FIC_2_APB_M_PRDATA[19]  (.D(\prdata[19] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[19]));
    SLE \pwdata[29]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[29]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[29]));
    SLE \paddr[5]  (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]), 
        .CLK(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d)
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_3));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[11]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[11]_net_1 ), .Y(\prdata[11] ));
    CFG3 #( .INIT(8'hA8) )  \prdata_0_iv_0_a2_0_0[16]  (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .C(
        CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET), .Y(
        \prdata_0_iv_0_a2_0[16] ));
    CFG4 #( .INIT(16'h0100) )  MDDR_PSEL_0_a4 (.A(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_10), .C(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11), .D(psel_net_1), .Y(
        CORECONFIGP_0_MDDR_APBmslave_PSELx));
    SLE \paddr[2]  (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), 
        .CLK(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d)
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_0));
    CFG2 #( .INIT(4'h8) )  \prdata_0_iv_0_a2_0[1]  (.A(N_126), .B(
        CORECONFIGP_0_SOFT_RESET_F2M), .Y(N_115));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[7]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[7]), .B(
        CORECONFIGP_0_SOFT_SDIF0_PHY_RESET), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[7]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[13]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[13]), .B(
        \soft_reset_reg[13]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[13]_net_1 ));
    SLE \pwdata[24]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[24]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[24]));
    SLE \FIC_2_APB_M_PRDATA[26]  (.D(\prdata[26] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[26]));
    SLE \FIC_2_APB_M_PRDATA[21]  (.D(\prdata[21] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[21]));
    CFG2 #( .INIT(4'h4) )  soft_reset_reg6_0_a2_0 (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .Y(
        soft_reset_reg6_0_a2_0_net_1));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[25]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[25]), .Y(\prdata[25] ));
    CFG2 #( .INIT(4'hE) )  state_s0_0_a2_0_a2_i (.A(\state[1]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(state_347_d_i_0));
    SLE \control_reg_1[1]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(control_reg_15), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(CORECONFIGP_0_CONFIG2_DONE)
        );
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[6]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[6]_net_1 ), .Y(\prdata[6] ));
    SLE \FIC_2_APB_M_PRDATA[22]  (.D(\prdata[22] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[22]));
    SLE FIC_2_APB_M_PREADY (.D(\state[1]_net_1 ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(N_51_i_0), .ALn(
        MSS_ADLIB_INST_RNI7K43), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY));
    SLE \pwdata[8]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[8]));
    SLE \FIC_2_APB_M_PRDATA[20]  (.D(\prdata[20] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[20]));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[0]  (.A(
        \prdata_0_iv_0_tz[0]_net_1 ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[0]), .C(N_39), .D(N_38), .Y(
        \prdata_0_iv_0_0[0]_net_1 ));
    CFG4 #( .INIT(16'h8F88) )  psel_RNIPEDQ (.A(psel_net_1), .B(
        g1_0_0_0), .C(CORECONFIGP_0_MDDR_APBmslave_PREADY), .D(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .Y(N_46));
    CFG4 #( .INIT(16'hF888) )  pslverr_0_iv_0_0 (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR), .B(N_39), .C(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .D(
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR), .Y(pslverr));
    CFG4 #( .INIT(16'h0010) )  \prdata_0_iv_0_a2_1_s[0]  (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .C(
        CORECONFIGP_0_CONFIG1_DONE), .D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]), .Y(
        prdata_0_iv_0_a2_1_out));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[6]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[6]), .B(
        \soft_reset_reg[6]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[6]_net_1 ));
    SLE \FIC_2_APB_M_PRDATA[23]  (.D(\prdata[23] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[23]));
    GND GND (.Y(GND_net_1));
    SLE \FIC_2_APB_M_PRDATA[17]  (.D(\prdata[17] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]));
    SLE \pwdata[10]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[10]));
    SLE \FIC_2_APB_M_PRDATA[29]  (.D(\prdata[29] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[29]));
    CFG3 #( .INIT(8'h40) )  \prdata_0_iv_0_a2_1_0[5]  (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]), .C(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .Y(
        \prdata_0_iv_0_a2_1[5] ));
    SLE \pwdata[4]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[4]));
    CFG3 #( .INIT(8'h04) )  \prdata_0_iv_0_a3_s_0[2]  (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .C(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]), .Y(
        prdata_0_iv_0_a3_out_0));
    CFG2 #( .INIT(4'h8) )  \prdata_0_iv_0_a2_2[5]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .Y(N_113));
    SLE \soft_reset_reg[6]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[6]_net_1 ));
    SLE \pwdata[7]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[7]));
    SLE MDDR_PENABLE (.D(MDDR_PENABLE_2), .CLK(un1_M2S_MSS_sb_0_4_i_0), 
        .EN(VCC_net_1), .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CORECONFIGP_0_MDDR_APBmslave_PENABLE));
    SLE \paddr[7]  (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]), 
        .CLK(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d)
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_5));
    SLE \pwdata[0]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[0]));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[7]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[7]_net_1 ), .Y(\prdata[7] ));
    SLE \pwdata[13]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[13]));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[20]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[20]), .Y(\prdata[20] ));
    SLE \soft_reset_reg[3]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[3]_net_1 ));
    SLE \soft_reset_reg[15]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET));
    SLE SDIF0_PENABLE (.D(N_16_i_0), .CLK(un1_M2S_MSS_sb_0_4_i_0), .EN(
        VCC_net_1), .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE));
    SLE \paddr[12]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_10));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[26]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[26]), .Y(\prdata[26] ));
    SLE \pwdata[30]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[30]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[30]));
    SLE \FIC_2_APB_M_PRDATA[31]  (.D(\prdata[31] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[31]));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[22]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[22]), .Y(\prdata[22] ));
    SLE psel (.D(state_347_d_i_0), .CLK(un1_M2S_MSS_sb_0_4_i_0), .EN(
        VCC_net_1), .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        psel_net_1));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[23]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[23]), .Y(\prdata[23] ));
    SLE \soft_reset_reg[2]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CORECONFIGP_0_SOFT_M3_RESET));
    CFG3 #( .INIT(8'h53) )  FIC_2_APB_M_PREADY_RNO (.A(N_46), .B(N_50), 
        .C(\state[1]_net_1 ), .Y(N_51_i_0));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[14]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[14]), .B(
        \soft_reset_reg[14]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[14]_net_1 ));
    SLE \paddr[13]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11));
    SLE \pwdata[20]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[20]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[20]));
    CFG4 #( .INIT(16'h0100) )  MDDR_PENABLE_2_0_a2 (.A(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_10), .C(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11), .D(\state[1]_net_1 ), 
        .Y(MDDR_PENABLE_2));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[9]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[9]), .B(
        \soft_reset_reg[9]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[9]_net_1 ));
    SLE \FIC_2_APB_M_PRDATA[18]  (.D(\prdata[18] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[18]));
    SLE \pwdata[17]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[17]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[17]));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[15]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[15]_net_1 ), .Y(\prdata[15] ));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0[18]  (.A(
        \prdata_0_iv_0_a2_0[17] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[18]), .C(N_39), .D(N_122), 
        .Y(\prdata[18] ));
    SLE \soft_reset_reg[14]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[14]_net_1 )
        );
    SLE \FIC_2_APB_M_PRDATA[30]  (.D(\prdata[30] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[30]));
    CFG1 #( .INIT(2'h1) )  \soft_reset_reg_RNI6AJD[2]  (.A(
        CORECONFIGP_0_SOFT_M3_RESET), .Y(
        CORECONFIGP_0_SOFT_M3_RESET_i_0));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[10]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[10]_net_1 ), .Y(\prdata[10] ));
    SLE \pwdata[23]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[23]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[23]));
    CFG4 #( .INIT(16'h30B0) )  \prdata_0_iv_0_a3[2]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11), .B(psel_net_1), .C(
        prdata_0_iv_0_a3_out_0), .D(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .Y(N_126));
    SLE \soft_reset_reg[8]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[8]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[21]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[21]), .Y(\prdata[21] ));
    SLE \FIC_2_APB_M_PRDATA[27]  (.D(\prdata[27] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[27]));
    SLE \FIC_2_APB_M_PRDATA[4]  (.D(\prdata[4] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[4]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[4]), .B(
        \soft_reset_reg[4]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[4]_net_1 ));
    SLE \soft_reset_reg[0]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[3]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[3]_net_1 ), .Y(\prdata[3] ));
    SLE \pwdata[27]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[27]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[27]));
    CFG4 #( .INIT(16'hFFF8) )  \prdata_0_iv_0[5]  (.A(
        \soft_reset_reg[5]_net_1 ), .B(N_126), .C(
        \prdata_0_iv_0_0[5]_net_1 ), .D(N_113), .Y(\prdata[5] ));
    SLE \pwdata[1]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[1]));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[9]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[9]_net_1 ), .Y(\prdata[9] ));
    CFG3 #( .INIT(8'h4F) )  \prdata_0_iv_0_o4[0]  (.A(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11), .C(psel_net_1), .Y(N_38)
        );
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0[17]  (.A(
        \prdata_0_iv_0_a2_0[17] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[17]), .C(N_39), .D(N_122), 
        .Y(\prdata[17] ));
    SLE \soft_reset_reg[1]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CORECONFIGP_0_SOFT_RESET_F2M));
    SLE \paddr[9]  (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]), 
        .CLK(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d)
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_7));
    SLE \FIC_2_APB_M_PRDATA[28]  (.D(\prdata[28] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[28]));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[1]  (.A(
        \prdata_0_iv_0_a2_1[1] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[1]), .C(N_39), .D(N_38), .Y(
        \prdata_0_iv_0_0[1]_net_1 ));
    SLE \paddr[15]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ));
    SLE \pwdata[16]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[16]));
    SLE \FIC_2_APB_M_PRDATA[3]  (.D(\prdata[3] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]));
    SLE \FIC_2_APB_M_PRDATA[14]  (.D(\prdata[14] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[2]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[2]_net_1 ), .Y(\prdata[2] ));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[4]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[4]_net_1 ), .Y(\prdata[4] ));
    CFG3 #( .INIT(8'hFD) )  \state_RNIOPSK[0]  (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE), .C(
        \state[0]_net_1 ), .Y(N_50));
    SLE \paddr[11]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[11]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_9));
    SLE \control_reg_1[0]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(control_reg_15), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(CORECONFIGP_0_CONFIG1_DONE)
        );
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[10]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[10]), .B(
        \soft_reset_reg[10]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[10]_net_1 ));
    SLE \soft_reset_reg[5]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[5]_net_1 ));
    SLE \FIC_2_APB_M_PRDATA[15]  (.D(\prdata[15] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]));
    SLE \paddr[3]  (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]), 
        .CLK(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d)
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_1));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[19]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[19]), .Y(\prdata[19] ));
    SLE INIT_DONE_q2 (.D(INIT_DONE_q1_net_1), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(VCC_net_1), .ALn(
        MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INIT_DONE_q2_net_1));
    SLE pwrite (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE));
    CFG4 #( .INIT(16'h5040) )  \prdata_0_iv_0_a2_1[0]  (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]), .C(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .D(
        INIT_DONE_q2_net_1), .Y(\prdata_0_iv_0_a2_1[0]_net_1 ));
    SLE \soft_reset_reg[10]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[10]_net_1 )
        );
    SLE \soft_reset_reg[4]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[4]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[12]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[12]), .B(
        \soft_reset_reg[12]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[12]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[13]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[13]_net_1 ), .Y(\prdata[13] ));
    SLE \FIC_2_APB_M_PRDATA[7]  (.D(\prdata[7] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]));
    SLE SDIF_RELEASED_q1 (.D(CORERESETP_0_SDIF_RELEASED), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(VCC_net_1), .ALn(
        MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(SDIF_RELEASED_q1_net_1));
    SLE \pwdata[26]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[26]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[26]));
    SLE \pwdata[6]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[6]));
    CFG4 #( .INIT(16'hFEFC) )  \prdata_0_iv_0[1]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .B(N_115), .C(
        \prdata_0_iv_0_0[1]_net_1 ), .D(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]), .Y(\prdata[1] ));
    SLE \pwdata[18]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[18]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[18]));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[12]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[12]_net_1 ), .Y(\prdata[12] ));
    SLE \pwdata[11]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[11]));
    SLE \paddr[6]  (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]), 
        .CLK(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d)
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_4));
    SLE \pwdata[12]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[12]));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv[0]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[0]_net_1 ), .Y(\prdata[0] ));
    CFG4 #( .INIT(16'h0080) )  control_reg_15_0_a2 (.A(
        control_reg_15_4), .B(psel_net_1), .C(
        control_reg_15_0_a2_0_net_1), .D(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .Y(control_reg_15));
    SLE \paddr[4]  (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), 
        .CLK(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d)
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_2));
    SLE \FIC_2_APB_M_PRDATA[24]  (.D(\prdata[24] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[24]));
    CFG4 #( .INIT(16'hECA0) )  \prdata_0_iv_0_0[5]  (.A(
        \prdata_0_iv_0_a2_1[5] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[5]), .C(N_38), .D(N_39), .Y(
        \prdata_0_iv_0_0[5]_net_1 ));
    SLE \FIC_2_APB_M_PRDATA[9]  (.D(\prdata[9] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]));
    CFG3 #( .INIT(8'hE2) )  \prdata_0_iv_0_m4[1]  (.A(
        CORECONFIGP_0_CONFIG2_DONE), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .C(
        SDIF_RELEASED_q2_net_1), .Y(N_48));
    SLE \pwdata[9]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[9]));
    CFG3 #( .INIT(8'hEA) )  \state_ns_0_0[1]  (.A(\state[0]_net_1 ), 
        .B(\state[1]_net_1 ), .C(N_46), .Y(\state_ns[1] ));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[29]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[29]), .Y(\prdata[29] ));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[28]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[28]), .Y(\prdata[28] ));
    SLE \state[1]  (.D(\state_ns[1] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(VCC_net_1), .ALn(
        MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\state[1]_net_1 ));
    SLE \soft_reset_reg[13]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[13]_net_1 )
        );
    SLE \FIC_2_APB_M_PRDATA[25]  (.D(\prdata[25] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[25]));
    SLE \FIC_2_APB_M_PRDATA[1]  (.D(\prdata[1] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]));
    SLE \pwdata[31]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[31]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[31]));
    SLE \pwdata[28]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[28]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[28]));
    SLE \pwdata[15]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[15]));
    CFG4 #( .INIT(16'hECA0) )  \prdata_0_iv_0[16]  (.A(
        \prdata_0_iv_0_a2_0[16] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[16]), .C(N_122), .D(N_39), 
        .Y(\prdata[16] ));
    SLE \pwdata[5]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[5]));
    SLE INIT_DONE_q1 (.D(INIT_DONE_int), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(VCC_net_1), .ALn(
        MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INIT_DONE_q1_net_1));
    SLE \FIC_2_APB_M_PRDATA[8]  (.D(\prdata[8] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]));
    CFG2 #( .INIT(4'h8) )  R_SDIF0_PSEL_1_i_o2 (.A(psel_net_1), .B(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .Y(N_39));
    SLE \FIC_2_APB_M_PRDATA[5]  (.D(\prdata[5] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]));
    SLE \pwdata[21]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[21]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[21]));
    SLE \pwdata[22]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[22]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[22]));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[2]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[2]), .B(
        CORECONFIGP_0_SOFT_M3_RESET), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[2]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \paddr_RNIVFTE[15]  (.A(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY), .Y(g1_0_0_0));
    CFG2 #( .INIT(4'h1) )  
        un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_a3_0_a2 (.A(
        \state[1]_net_1 ), .B(N_50), .Y(\state_ns[0] ));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[30]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[30]), .Y(\prdata[30] ));
    CFG2 #( .INIT(4'h8) )  \prdata_0_iv_0_a2_0_0[17]  (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .Y(
        \prdata_0_iv_0_a2_0[17] ));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[15]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[15]), .B(
        CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET), .C(N_126), .D(N_39), 
        .Y(\prdata_0_iv_0_0[15]_net_1 ));
    SLE \FIC_2_APB_M_PRDATA[0]  (.D(\prdata[0] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]));
    CFG3 #( .INIT(8'hEC) )  \prdata_0_iv_0[8]  (.A(N_126), .B(
        \prdata_0_iv_0_0[8]_net_1 ), .C(\soft_reset_reg[8]_net_1 ), .Y(
        \prdata[8] ));
    SLE \paddr[14]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[14]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_12));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[24]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[24]), .Y(\prdata[24] ));
    CFG4 #( .INIT(16'h4000) )  control_reg_15_0_a2_4 (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11), .C(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE), .D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE), .Y(
        control_reg_15_4));
    SLE \FIC_2_APB_M_PRDATA[16]  (.D(\prdata[16] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]));
    SLE \paddr[10]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_8));
    SLE \FIC_2_APB_M_PRDATA[11]  (.D(\prdata[11] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]));
    CFG2 #( .INIT(4'h2) )  \prdata_0_iv_0_a3_0[0]  (.A(N_38), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]), .Y(N_122));
    CFG4 #( .INIT(16'hF888) )  \prdata_0_iv_0_0[8]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[8]), .C(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]), .D(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .Y(
        \prdata_0_iv_0_0[8]_net_1 ));
    SLE \soft_reset_reg[9]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[9]_net_1 ));
    SLE \soft_reset_reg[11]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[11]_net_1 )
        );
    SLE \pwdata[2]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[2]));
    SLE \FIC_2_APB_M_PRDATA[6]  (.D(\prdata[6] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]));
    SLE \pwdata[19]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[19]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[19]));
    SLE \pwdata[25]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[25]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[25]));
    SLE \FIC_2_APB_M_PRDATA[2]  (.D(\prdata[2] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]));
    SLE \soft_reset_reg[16]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET));
    CFG3 #( .INIT(8'hF8) )  \prdata_0_iv_0[14]  (.A(
        CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]), .B(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .C(
        \prdata_0_iv_0_0[14]_net_1 ), .Y(\prdata[14] ));
    SLE \pwdata[14]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[14]));
    SLE \FIC_2_APB_M_PRDATA[12]  (.D(\prdata[12] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]));
    SLE SDIF_RELEASED_q2 (.D(SDIF_RELEASED_q1_net_1), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(VCC_net_1), .ALn(
        MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(SDIF_RELEASED_q2_net_1));
    CFG3 #( .INIT(8'h04) )  \prdata_0_iv_0_a2_1_0[1]  (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]), .B(N_48), .C(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .Y(
        \prdata_0_iv_0_a2_1[1] ));
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[3]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[3]), .B(
        \soft_reset_reg[3]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[3]_net_1 ));
    CFG2 #( .INIT(4'h1) )  state_s0_0_a2_0_a2 (.A(\state[1]_net_1 ), 
        .B(\state[0]_net_1 ), .Y(state_347_d));
    CFG4 #( .INIT(16'h2000) )  soft_reset_reg6_0_a2 (.A(
        soft_reset_reg6_0_a2_0_net_1), .B(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .C(control_reg_15_4), 
        .D(psel_net_1), .Y(soft_reset_reg6));
    SLE \FIC_2_APB_M_PRDATA[10]  (.D(\prdata[10] ), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]));
    SLE \pwdata[3]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[3]));
    CFG1 #( .INIT(2'h1) )  \soft_reset_reg_RNI59JD[1]  (.A(
        CORECONFIGP_0_SOFT_RESET_F2M), .Y(
        CORECONFIGP_0_SOFT_RESET_F2M_i_0));
    SLE \paddr[8]  (.D(M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]), 
        .CLK(FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(state_347_d)
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_6));
    CFG2 #( .INIT(4'h8) )  \FIC_2_APB_M_PRDATA_RNO[31]  (.A(N_39), .B(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[31]), .Y(\prdata[31] ));
    SLE \soft_reset_reg[7]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CORECONFIGP_0_SOFT_SDIF0_PHY_RESET));
    SLE \soft_reset_reg[12]  (.D(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(soft_reset_reg6), 
        .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\soft_reset_reg[12]_net_1 )
        );
    CFG4 #( .INIT(16'hEAC0) )  \prdata_0_iv_0_0[11]  (.A(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[11]), .B(
        \soft_reset_reg[11]_net_1 ), .C(N_126), .D(N_39), .Y(
        \prdata_0_iv_0_0[11]_net_1 ));
    CFG2 #( .INIT(4'h1) )  control_reg_15_0_a2_0 (.A(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]), .B(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]), .Y(
        control_reg_15_0_a2_0_net_1));
    SLE FIC_2_APB_M_PSLVERR (.D(pslverr), .CLK(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), .EN(\state[1]_net_1 )
        , .ALn(MSS_ADLIB_INST_RNI7K43), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR));
    CFG2 #( .INIT(4'h8) )  SDIF0_PENABLE_RNO (.A(\state[1]_net_1 ), .B(
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[15] ), .Y(N_16_i_0));
    
endmodule


module M2S_MSS_sb(
       M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA,
       MDDR_DQ,
       MDDR_DM_RDQS,
       MDDR_BA,
       MDDR_ADDR,
       MDDR_DQS_N,
       MDDR_DQS,
       DEVRST_N,
       FAB_CCC_GL0_c,
       FAB_CCC_LOCK_c,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY,
       N_39,
       M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR,
       SDIF0_SPLL_LOCK_c,
       SDIF0_1_CORE_RESET_N_c,
       SDIF0_0_CORE_RESET_N_c,
       SDIF0_PHY_RESET_N_c,
       SPI_1_SS0,
       SPI_1_DO,
       SPI_1_DI,
       SPI_1_CLK,
       SPI_0_SS0,
       SPI_0_DO,
       SPI_0_DI,
       SPI_0_CLK,
       MMUART_1_TXD,
       MMUART_1_RXD,
       MMUART_0_TXD,
       MMUART_0_RXD,
       MDDR_WE_N,
       MDDR_RESET_N,
       MDDR_RAS_N,
       MDDR_ODT,
       MDDR_DQS_TMATCH_0_OUT,
       MDDR_DQS_TMATCH_0_IN,
       MDDR_CS_N,
       MDDR_CKE,
       MDDR_CAS_N,
       I2C_1_SDA,
       I2C_1_SCL,
       I2C_0_SDA,
       I2C_0_SCL,
       GPIO_3_M2F_c,
       GPIO_2_M2F_c,
       GPIO_1_M2F_c,
       GPIO_0_M2F_c,
       MDDR_CLK_N,
       MDDR_CLK
    );
output [14:2] M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR;
output [31:0] M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA;
input  [31:0] M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA;
inout  [7:0] MDDR_DQ;
inout  [0:0] MDDR_DM_RDQS;
output [2:0] MDDR_BA;
output [15:0] MDDR_ADDR;
inout  [0:0] MDDR_DQS_N;
inout  [0:0] MDDR_DQS;
input  DEVRST_N;
output FAB_CCC_GL0_c;
inout  FAB_CCC_LOCK_c;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE;
output M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE;
input  M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY;
output N_39;
input  M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR;
input  SDIF0_SPLL_LOCK_c;
output SDIF0_1_CORE_RESET_N_c;
output SDIF0_0_CORE_RESET_N_c;
output SDIF0_PHY_RESET_N_c;
inout  SPI_1_SS0;
output SPI_1_DO;
input  SPI_1_DI;
inout  SPI_1_CLK;
inout  SPI_0_SS0;
output SPI_0_DO;
input  SPI_0_DI;
inout  SPI_0_CLK;
output MMUART_1_TXD;
input  MMUART_1_RXD;
output MMUART_0_TXD;
input  MMUART_0_RXD;
output MDDR_WE_N;
output MDDR_RESET_N;
output MDDR_RAS_N;
output MDDR_ODT;
output MDDR_DQS_TMATCH_0_OUT;
input  MDDR_DQS_TMATCH_0_IN;
output MDDR_CS_N;
output MDDR_CKE;
output MDDR_CAS_N;
inout  I2C_1_SDA;
inout  I2C_1_SCL;
inout  I2C_0_SDA;
inout  I2C_0_SCL;
output GPIO_3_M2F_c;
output GPIO_2_M2F_c;
output GPIO_1_M2F_c;
output GPIO_0_M2F_c;
output MDDR_CLK_N;
output MDDR_CLK;

    wire SYSRESET_POR_net_1, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[17] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[18] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[19] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[20] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[21] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[22] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[23] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[24] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[25] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[26] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[27] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[28] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[29] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[30] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[31] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[18] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[19] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[20] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[21] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[22] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[23] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[24] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[25] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[26] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[27] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[28] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[29] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[30] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[31] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15] , 
        CORECONFIGP_0_SOFT_RESET_F2M_i_0, 
        CORECONFIGP_0_SOFT_M3_RESET_i_0, MSS_ADLIB_INST_RNI7K43, 
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA, 
        CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET, 
        CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET, 
        CORECONFIGP_0_CONFIG1_DONE, CORECONFIGP_0_CONFIG2_DONE, 
        CORECONFIGP_0_SOFT_SDIF0_PHY_RESET, 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        un1_M2S_MSS_sb_0_4_i_0, INIT_DONE_int, 
        CORERESETP_0_SDIF_RELEASED, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        FABOSC_0_RCOSC_25_50MHZ_O2F, 
        M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F, GND_net_1, VCC_net_1;
    
    M2S_MSS_sb_FABOSC_0_OSC FABOSC_0 (.FABOSC_0_RCOSC_25_50MHZ_O2F(
        FABOSC_0_RCOSC_25_50MHZ_O2F), 
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    CoreResetP_Z2 CORERESETP_0 (.FAB_CCC_GL0_c(FAB_CCC_GL0_c), 
        .CORERESETP_0_SDIF_RELEASED(CORERESETP_0_SDIF_RELEASED), 
        .FABOSC_0_RCOSC_25_50MHZ_O2F(FABOSC_0_RCOSC_25_50MHZ_O2F), 
        .INIT_DONE_int(INIT_DONE_int), .SYSRESET_POR(
        SYSRESET_POR_net_1), .M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F(
        M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F), .MSS_ADLIB_INST_RNI7K43(
        MSS_ADLIB_INST_RNI7K43), .CORECONFIGP_0_CONFIG1_DONE(
        CORECONFIGP_0_CONFIG1_DONE), .CORECONFIGP_0_CONFIG2_DONE(
        CORECONFIGP_0_CONFIG2_DONE), .SDIF0_SPLL_LOCK_c(
        SDIF0_SPLL_LOCK_c), .CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET(
        CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET), 
        .SDIF0_1_CORE_RESET_N_c(SDIF0_1_CORE_RESET_N_c), 
        .CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET(
        CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET), 
        .SDIF0_0_CORE_RESET_N_c(SDIF0_0_CORE_RESET_N_c), 
        .CORECONFIGP_0_SOFT_SDIF0_PHY_RESET(
        CORECONFIGP_0_SOFT_SDIF0_PHY_RESET), .SDIF0_PHY_RESET_N_c(
        SDIF0_PHY_RESET_N_c));
    VCC VCC (.Y(VCC_net_1));
    M2S_MSS_sb_MSS M2S_MSS_sb_MSS_0 (.MDDR_DQ({MDDR_DQ[7], MDDR_DQ[6], 
        MDDR_DQ[5], MDDR_DQ[4], MDDR_DQ[3], MDDR_DQ[2], MDDR_DQ[1], 
        MDDR_DQ[0]}), .MDDR_DM_RDQS({MDDR_DM_RDQS[0]}), .MDDR_BA({
        MDDR_BA[2], MDDR_BA[1], MDDR_BA[0]}), .MDDR_ADDR({
        MDDR_ADDR[15], MDDR_ADDR[14], MDDR_ADDR[13], MDDR_ADDR[12], 
        MDDR_ADDR[11], MDDR_ADDR[10], MDDR_ADDR[9], MDDR_ADDR[8], 
        MDDR_ADDR[7], MDDR_ADDR[6], MDDR_ADDR[5], MDDR_ADDR[4], 
        MDDR_ADDR[3], MDDR_ADDR[2], MDDR_ADDR[1], MDDR_ADDR[0]}), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR({
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2] }), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA({
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[31] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[30] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[29] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[28] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[27] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[26] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[25] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[24] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[23] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[22] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[21] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[20] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[19] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[18] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[17] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0] }), 
        .CORECONFIGP_0_MDDR_APBmslave_PRDATA({
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0] }), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA({
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[31] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[30] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[29] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[28] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[27] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[26] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[25] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[24] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[23] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[22] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[21] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[20] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[19] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[18] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR({
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[2]}), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA({
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[15], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[14], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[13], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[12], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[11], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[2], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[1], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[0]}), .MDDR_DQS_N({
        MDDR_DQS_N[0]}), .MDDR_DQS({MDDR_DQS[0]}), 
        .FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), 
        .MSS_ADLIB_INST_RNI7K43(MSS_ADLIB_INST_RNI7K43), 
        .un1_M2S_MSS_sb_0_4_i_0(un1_M2S_MSS_sb_0_4_i_0), .SPI_1_SS0(
        SPI_1_SS0), .SPI_1_DO(SPI_1_DO), .SPI_1_DI(SPI_1_DI), 
        .SPI_1_CLK(SPI_1_CLK), .SPI_0_SS0(SPI_0_SS0), .SPI_0_DO(
        SPI_0_DO), .SPI_0_DI(SPI_0_DI), .SPI_0_CLK(SPI_0_CLK), 
        .MMUART_1_TXD(MMUART_1_TXD), .MMUART_1_RXD(MMUART_1_RXD), 
        .MMUART_0_TXD(MMUART_0_TXD), .MMUART_0_RXD(MMUART_0_RXD), 
        .MDDR_WE_N(MDDR_WE_N), .MDDR_RESET_N(MDDR_RESET_N), 
        .MDDR_RAS_N(MDDR_RAS_N), .MDDR_ODT(MDDR_ODT), 
        .MDDR_DQS_TMATCH_0_OUT(MDDR_DQS_TMATCH_0_OUT), 
        .MDDR_DQS_TMATCH_0_IN(MDDR_DQS_TMATCH_0_IN), .MDDR_CS_N(
        MDDR_CS_N), .MDDR_CKE(MDDR_CKE), .MDDR_CAS_N(MDDR_CAS_N), 
        .I2C_1_SDA(I2C_1_SDA), .I2C_1_SCL(I2C_1_SCL), .I2C_0_SDA(
        I2C_0_SDA), .I2C_0_SCL(I2C_0_SCL), .GPIO_3_M2F_c(GPIO_3_M2F_c), 
        .GPIO_2_M2F_c(GPIO_2_M2F_c), 
        .M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F(
        M2S_MSS_sb_MSS_TMP_0_MSS_RESET_N_M2F), .GPIO_1_M2F_c(
        GPIO_1_M2F_c), .GPIO_0_M2F_c(GPIO_0_M2F_c), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE), 
        .CORECONFIGP_0_MDDR_APBmslave_PREADY(
        CORECONFIGP_0_MDDR_APBmslave_PREADY), 
        .CORECONFIGP_0_MDDR_APBmslave_PSLVERR(
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR), 
        .CORECONFIGP_0_SOFT_M3_RESET_i_0(
        CORECONFIGP_0_SOFT_M3_RESET_i_0), .FAB_CCC_LOCK_c(
        FAB_CCC_LOCK_c), .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR), 
        .CORECONFIGP_0_SOFT_RESET_F2M_i_0(
        CORECONFIGP_0_SOFT_RESET_F2M_i_0), .FAB_CCC_GL0_c(
        FAB_CCC_GL0_c), .CORECONFIGP_0_MDDR_APBmslave_PENABLE(
        CORECONFIGP_0_MDDR_APBmslave_PENABLE), 
        .CORECONFIGP_0_MDDR_APBmslave_PSELx(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE), .MDDR_CLK_N(MDDR_CLK_N), 
        .MDDR_CLK(MDDR_CLK));
    M2S_MSS_sb_CCC_0_FCCC CCC_0 (.FAB_CCC_GL0_c(FAB_CCC_GL0_c), 
        .FAB_CCC_LOCK_c(FAB_CCC_LOCK_c), 
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    GND GND (.Y(GND_net_1));
    CoreConfigP_Z1 CORECONFIGP_0 (
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR({
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA({
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[31], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[30], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[29], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[28], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[27], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[26], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[25], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[24], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[23], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[22], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[21], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[20], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[19], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[18], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[17], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[16], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[15], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[14], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[13], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[12], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[11], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[2], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[1], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[0]}), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA({
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[31] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[30] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[29] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[28] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[27] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[26] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[25] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[24] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[23] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[22] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[21] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[20] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[19] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[18] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[17] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0] }), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA({
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[31] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[30] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[29] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[28] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[27] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[26] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[25] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[24] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[23] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[22] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[21] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[20] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[19] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[18] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1] , 
        \M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA({
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[31], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[30], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[29], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[28], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[27], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[26], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[25], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[24], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[23], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[22], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[21], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[20], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[19], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[18], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[17], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[16], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[15], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[14], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[13], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[12], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[11], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[10], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[9], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[8], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[7], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[6], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[5], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[4], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[3], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[2], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[1], 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[0]}), 
        .CORECONFIGP_0_MDDR_APBmslave_PRDATA({
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1] , 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_6(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[8]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_7(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[9]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_8(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[10]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_9(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[11]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_10(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[12]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_11(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[13]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_12(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[14]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_0(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[2]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_1(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[3]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_2(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[4]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_3(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[5]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_4(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[6]), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR_5(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[7]), 
        .CORECONFIGP_0_SOFT_RESET_F2M_i_0(
        CORECONFIGP_0_SOFT_RESET_F2M_i_0), 
        .CORECONFIGP_0_SOFT_M3_RESET_i_0(
        CORECONFIGP_0_SOFT_M3_RESET_i_0), .MSS_ADLIB_INST_RNI7K43(
        MSS_ADLIB_INST_RNI7K43), 
        .FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA(
        FIC_2_APB_M_PCLK_inferred_clock_RNIVUHA), 
        .CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET(
        CORECONFIGP_0_SOFT_SDIF0_0_CORE_RESET), 
        .CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET(
        CORECONFIGP_0_SOFT_SDIF0_1_CORE_RESET), 
        .CORECONFIGP_0_CONFIG1_DONE(CORECONFIGP_0_CONFIG1_DONE), 
        .CORECONFIGP_0_CONFIG2_DONE(CORECONFIGP_0_CONFIG2_DONE), 
        .CORECONFIGP_0_SOFT_SDIF0_PHY_RESET(
        CORECONFIGP_0_SOFT_SDIF0_PHY_RESET), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE), 
        .un1_M2S_MSS_sb_0_4_i_0(un1_M2S_MSS_sb_0_4_i_0), 
        .INIT_DONE_int(INIT_DONE_int), .CORERESETP_0_SDIF_RELEASED(
        CORERESETP_0_SDIF_RELEASED), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE), 
        .CORECONFIGP_0_MDDR_APBmslave_PENABLE(
        CORECONFIGP_0_MDDR_APBmslave_PENABLE), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx), 
        .M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE(
        M2S_MSS_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE), 
        .CORECONFIGP_0_MDDR_APBmslave_PREADY(
        CORECONFIGP_0_MDDR_APBmslave_PREADY), 
        .CORECONFIGP_0_MDDR_APBmslave_PSELx(
        CORECONFIGP_0_MDDR_APBmslave_PSELx), .N_39(N_39), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR), 
        .CORECONFIGP_0_MDDR_APBmslave_PSLVERR(
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR));
    SYSRESET SYSRESET_POR (.POWER_ON_RESET_N(SYSRESET_POR_net_1), 
        .DEVRST_N(DEVRST_N));
    
endmodule


module M2S_MSS(
       PCIE_0_INTERRUPT,
       MDDR_ADDR,
       MDDR_BA,
       MDDR_DM_RDQS,
       MDDR_DQ,
       MDDR_DQS,
       MDDR_DQS_N,
       APB_S_PCLK,
       APB_S_PRESET_N,
       CLK_BASE,
       DEVRST_N,
       MDDR_DQS_TMATCH_0_IN,
       MMUART_0_RXD,
       MMUART_1_RXD,
       PCIE_0_CORE_RESET_N,
       PCIE_0_PERST_N,
       PHY_RESET_N,
       REFCLK0_N,
       REFCLK0_P,
       RXD0_N,
       RXD0_P,
       RXD1_N,
       RXD1_P,
       RXD2_N,
       RXD2_P,
       RXD3_N,
       RXD3_P,
       SDIF0_SPLL_LOCK,
       SPI_0_DI,
       SPI_1_DI,
       FAB_CCC_GL0,
       FAB_CCC_LOCK,
       GPIO_0_M2F,
       GPIO_1_M2F,
       GPIO_2_M2F,
       GPIO_3_M2F,
       MDDR_CAS_N,
       MDDR_CKE,
       MDDR_CLK,
       MDDR_CLK_N,
       MDDR_CS_N,
       MDDR_DQS_TMATCH_0_OUT,
       MDDR_ODT,
       MDDR_RAS_N,
       MDDR_RESET_N,
       MDDR_WE_N,
       MMUART_0_TXD,
       MMUART_1_TXD,
       SDIF0_0_CORE_RESET_N,
       SDIF0_1_CORE_RESET_N,
       SDIF0_PHY_RESET_N,
       SPI_0_DO,
       SPI_1_DO,
       TXD0_N,
       TXD0_P,
       TXD1_N,
       TXD1_P,
       TXD2_N,
       TXD2_P,
       TXD3_N,
       TXD3_P,
       I2C_0_SCL,
       I2C_0_SDA,
       I2C_1_SCL,
       I2C_1_SDA,
       SPI_0_CLK,
       SPI_0_SS0,
       SPI_1_CLK,
       SPI_1_SS0
    );
input  [3:0] PCIE_0_INTERRUPT;
output [15:0] MDDR_ADDR;
output [2:0] MDDR_BA;
inout  [0:0] MDDR_DM_RDQS;
inout  [7:0] MDDR_DQ;
inout  [0:0] MDDR_DQS;
inout  [0:0] MDDR_DQS_N;
input  APB_S_PCLK;
input  APB_S_PRESET_N;
input  CLK_BASE;
input  DEVRST_N;
input  MDDR_DQS_TMATCH_0_IN;
input  MMUART_0_RXD;
input  MMUART_1_RXD;
input  PCIE_0_CORE_RESET_N;
input  PCIE_0_PERST_N;
input  PHY_RESET_N;
input  REFCLK0_N;
input  REFCLK0_P;
input  RXD0_N;
input  RXD0_P;
input  RXD1_N;
input  RXD1_P;
input  RXD2_N;
input  RXD2_P;
input  RXD3_N;
input  RXD3_P;
input  SDIF0_SPLL_LOCK;
input  SPI_0_DI;
input  SPI_1_DI;
output FAB_CCC_GL0;
output FAB_CCC_LOCK;
output GPIO_0_M2F;
output GPIO_1_M2F;
output GPIO_2_M2F;
output GPIO_3_M2F;
output MDDR_CAS_N;
output MDDR_CKE;
output MDDR_CLK;
output MDDR_CLK_N;
output MDDR_CS_N;
output MDDR_DQS_TMATCH_0_OUT;
output MDDR_ODT;
output MDDR_RAS_N;
output MDDR_RESET_N;
output MDDR_WE_N;
output MMUART_0_TXD;
output MMUART_1_TXD;
output SDIF0_0_CORE_RESET_N;
output SDIF0_1_CORE_RESET_N;
output SDIF0_PHY_RESET_N;
output SPI_0_DO;
output SPI_1_DO;
output TXD0_N;
output TXD0_P;
output TXD1_N;
output TXD1_P;
output TXD2_N;
output TXD2_P;
output TXD3_N;
output TXD3_P;
inout  I2C_0_SCL;
inout  I2C_0_SDA;
inout  I2C_1_SCL;
inout  I2C_1_SDA;
inout  SPI_0_CLK;
inout  SPI_0_SS0;
inout  SPI_1_CLK;
inout  SPI_1_SS0;

    wire \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[0] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[1] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[2] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[14] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[15] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[16] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[17] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[18] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[19] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[20] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[21] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[22] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[23] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[24] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[25] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[26] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[27] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[28] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[29] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[30] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[31] , 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY, 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR, 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[2] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[14] , 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE, 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[0] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[1] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[2] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[14] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[15] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[16] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[17] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[18] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[19] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[20] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[21] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[22] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[23] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[24] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[25] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[26] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[27] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[28] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[29] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[30] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[31] , 
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE, GND_net_1, VCC_net_1, N_39, 
        APB_S_PCLK_c, APB_S_PRESET_N_c, CLK_BASE_c, 
        PCIE_0_CORE_RESET_N_c, \PCIE_0_INTERRUPT_c[0] , 
        \PCIE_0_INTERRUPT_c[1] , \PCIE_0_INTERRUPT_c[2] , 
        \PCIE_0_INTERRUPT_c[3] , PCIE_0_PERST_N_c, PHY_RESET_N_c, 
        SDIF0_SPLL_LOCK_c, FAB_CCC_GL0_c, FAB_CCC_LOCK_c, GPIO_0_M2F_c, 
        GPIO_1_M2F_c, GPIO_2_M2F_c, GPIO_3_M2F_c, 
        SDIF0_0_CORE_RESET_N_c, SDIF0_1_CORE_RESET_N_c, 
        SDIF0_PHY_RESET_N_c;
    
    OUTBUF SDIF0_PHY_RESET_N_obuf (.D(SDIF0_PHY_RESET_N_c), .PAD(
        SDIF0_PHY_RESET_N));
    OUTBUF GPIO_1_M2F_obuf (.D(GPIO_1_M2F_c), .PAD(GPIO_1_M2F));
    INBUF CLK_BASE_ibuf (.PAD(CLK_BASE), .Y(CLK_BASE_c));
    OUTBUF GPIO_2_M2F_obuf (.D(GPIO_2_M2F_c), .PAD(GPIO_2_M2F));
    INBUF \PCIE_0_INTERRUPT_ibuf[3]  (.PAD(PCIE_0_INTERRUPT[3]), .Y(
        \PCIE_0_INTERRUPT_c[3] ));
    OUTBUF FAB_CCC_LOCK_obuf (.D(FAB_CCC_LOCK_c), .PAD(FAB_CCC_LOCK));
    M2S_MSS_SERDES_IF2_0_SERDES_IF2 SERDES_IF2_0 (
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA({
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[31] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[30] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[29] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[28] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[27] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[26] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[25] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[24] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[23] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[22] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[21] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[20] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[19] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[18] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[17] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[16] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[15] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[14] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[2] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[1] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[0] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR({
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[14] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[2] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA({
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[31] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[30] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[29] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[28] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[27] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[26] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[25] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[24] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[23] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[22] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[21] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[20] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[19] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[18] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[17] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[16] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[15] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[14] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[2] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[1] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[0] }), .PCIE_0_INTERRUPT_c({
        \PCIE_0_INTERRUPT_c[3] , \PCIE_0_INTERRUPT_c[2] , 
        \PCIE_0_INTERRUPT_c[1] , \PCIE_0_INTERRUPT_c[0] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR), .APB_S_PCLK_c(
        APB_S_PCLK_c), .M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE), .N_39(N_39), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE), .APB_S_PRESET_N_c(
        APB_S_PRESET_N_c), .CLK_BASE_c(CLK_BASE_c), .PCIE_0_PERST_N_c(
        PCIE_0_PERST_N_c), .PCIE_0_CORE_RESET_N_c(
        PCIE_0_CORE_RESET_N_c), .PHY_RESET_N_c(PHY_RESET_N_c), .RXD3_P(
        RXD3_P), .RXD2_P(RXD2_P), .RXD1_P(RXD1_P), .RXD0_P(RXD0_P), 
        .RXD3_N(RXD3_N), .RXD2_N(RXD2_N), .RXD1_N(RXD1_N), .RXD0_N(
        RXD0_N), .TXD3_P(TXD3_P), .TXD2_P(TXD2_P), .TXD1_P(TXD1_P), 
        .TXD0_P(TXD0_P), .TXD3_N(TXD3_N), .TXD2_N(TXD2_N), .TXD1_N(
        TXD1_N), .TXD0_N(TXD0_N), .REFCLK0_N(REFCLK0_N), .REFCLK0_P(
        REFCLK0_P));
    OUTBUF SDIF0_0_CORE_RESET_N_obuf (.D(SDIF0_0_CORE_RESET_N_c), .PAD(
        SDIF0_0_CORE_RESET_N));
    OUTBUF FAB_CCC_GL0_obuf (.D(FAB_CCC_GL0_c), .PAD(FAB_CCC_GL0));
    INBUF PCIE_0_PERST_N_ibuf (.PAD(PCIE_0_PERST_N), .Y(
        PCIE_0_PERST_N_c));
    GND GND (.Y(GND_net_1));
    M2S_MSS_sb M2S_MSS_sb_0 (.M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR({
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[14] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PADDR[2] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA({
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[31] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[30] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[29] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[28] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[27] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[26] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[25] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[24] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[23] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[22] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[21] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[20] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[19] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[18] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[17] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[16] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[15] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[14] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[2] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[1] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PWDATA[0] }), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA({
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[31] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[30] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[29] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[28] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[27] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[26] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[25] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[24] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[23] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[22] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[21] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[20] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[19] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[18] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[17] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[16] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[15] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[14] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[13] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[12] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[11] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[10] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[9] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[8] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[7] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[6] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[5] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[4] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[3] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[2] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[1] , 
        \M2S_MSS_sb_0_SDIF0_INIT_APB_PRDATA[0] }), .MDDR_DQ({
        MDDR_DQ[7], MDDR_DQ[6], MDDR_DQ[5], MDDR_DQ[4], MDDR_DQ[3], 
        MDDR_DQ[2], MDDR_DQ[1], MDDR_DQ[0]}), .MDDR_DM_RDQS({
        MDDR_DM_RDQS[0]}), .MDDR_BA({MDDR_BA[2], MDDR_BA[1], 
        MDDR_BA[0]}), .MDDR_ADDR({MDDR_ADDR[15], MDDR_ADDR[14], 
        MDDR_ADDR[13], MDDR_ADDR[12], MDDR_ADDR[11], MDDR_ADDR[10], 
        MDDR_ADDR[9], MDDR_ADDR[8], MDDR_ADDR[7], MDDR_ADDR[6], 
        MDDR_ADDR[5], MDDR_ADDR[4], MDDR_ADDR[3], MDDR_ADDR[2], 
        MDDR_ADDR[1], MDDR_ADDR[0]}), .MDDR_DQS_N({MDDR_DQS_N[0]}), 
        .MDDR_DQS({MDDR_DQS[0]}), .DEVRST_N(DEVRST_N), .FAB_CCC_GL0_c(
        FAB_CCC_GL0_c), .FAB_CCC_LOCK_c(FAB_CCC_LOCK_c), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PWRITE), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PENABLE), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PREADY), .N_39(N_39), 
        .M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR(
        M2S_MSS_sb_0_SDIF0_INIT_APB_PSLVERR), .SDIF0_SPLL_LOCK_c(
        SDIF0_SPLL_LOCK_c), .SDIF0_1_CORE_RESET_N_c(
        SDIF0_1_CORE_RESET_N_c), .SDIF0_0_CORE_RESET_N_c(
        SDIF0_0_CORE_RESET_N_c), .SDIF0_PHY_RESET_N_c(
        SDIF0_PHY_RESET_N_c), .SPI_1_SS0(SPI_1_SS0), .SPI_1_DO(
        SPI_1_DO), .SPI_1_DI(SPI_1_DI), .SPI_1_CLK(SPI_1_CLK), 
        .SPI_0_SS0(SPI_0_SS0), .SPI_0_DO(SPI_0_DO), .SPI_0_DI(SPI_0_DI)
        , .SPI_0_CLK(SPI_0_CLK), .MMUART_1_TXD(MMUART_1_TXD), 
        .MMUART_1_RXD(MMUART_1_RXD), .MMUART_0_TXD(MMUART_0_TXD), 
        .MMUART_0_RXD(MMUART_0_RXD), .MDDR_WE_N(MDDR_WE_N), 
        .MDDR_RESET_N(MDDR_RESET_N), .MDDR_RAS_N(MDDR_RAS_N), 
        .MDDR_ODT(MDDR_ODT), .MDDR_DQS_TMATCH_0_OUT(
        MDDR_DQS_TMATCH_0_OUT), .MDDR_DQS_TMATCH_0_IN(
        MDDR_DQS_TMATCH_0_IN), .MDDR_CS_N(MDDR_CS_N), .MDDR_CKE(
        MDDR_CKE), .MDDR_CAS_N(MDDR_CAS_N), .I2C_1_SDA(I2C_1_SDA), 
        .I2C_1_SCL(I2C_1_SCL), .I2C_0_SDA(I2C_0_SDA), .I2C_0_SCL(
        I2C_0_SCL), .GPIO_3_M2F_c(GPIO_3_M2F_c), .GPIO_2_M2F_c(
        GPIO_2_M2F_c), .GPIO_1_M2F_c(GPIO_1_M2F_c), .GPIO_0_M2F_c(
        GPIO_0_M2F_c), .MDDR_CLK_N(MDDR_CLK_N), .MDDR_CLK(MDDR_CLK));
    INBUF \PCIE_0_INTERRUPT_ibuf[1]  (.PAD(PCIE_0_INTERRUPT[1]), .Y(
        \PCIE_0_INTERRUPT_c[1] ));
    INBUF \PCIE_0_INTERRUPT_ibuf[2]  (.PAD(PCIE_0_INTERRUPT[2]), .Y(
        \PCIE_0_INTERRUPT_c[2] ));
    INBUF APB_S_PRESET_N_ibuf (.PAD(APB_S_PRESET_N), .Y(
        APB_S_PRESET_N_c));
    INBUF SDIF0_SPLL_LOCK_ibuf (.PAD(SDIF0_SPLL_LOCK), .Y(
        SDIF0_SPLL_LOCK_c));
    INBUF \PCIE_0_INTERRUPT_ibuf[0]  (.PAD(PCIE_0_INTERRUPT[0]), .Y(
        \PCIE_0_INTERRUPT_c[0] ));
    INBUF PCIE_0_CORE_RESET_N_ibuf (.PAD(PCIE_0_CORE_RESET_N), .Y(
        PCIE_0_CORE_RESET_N_c));
    OUTBUF GPIO_0_M2F_obuf (.D(GPIO_0_M2F_c), .PAD(GPIO_0_M2F));
    VCC VCC (.Y(VCC_net_1));
    OUTBUF GPIO_3_M2F_obuf (.D(GPIO_3_M2F_c), .PAD(GPIO_3_M2F));
    INBUF APB_S_PCLK_ibuf (.PAD(APB_S_PCLK), .Y(APB_S_PCLK_c));
    OUTBUF SDIF0_1_CORE_RESET_N_obuf (.D(SDIF0_1_CORE_RESET_N_c), .PAD(
        SDIF0_1_CORE_RESET_N));
    INBUF PHY_RESET_N_ibuf (.PAD(PHY_RESET_N), .Y(PHY_RESET_N_c));
    
endmodule
