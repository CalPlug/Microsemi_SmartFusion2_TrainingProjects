`timescale 1 ns/100 ps
// Version: 


module SERDESIF_075(
       APB_PRDATA,
       APB_PREADY,
       APB_PSLVERR,
       ATXCLKSTABLE,
       EPCS_READY,
       EPCS_RXCLK,
       EPCS_RXCLK_0,
       EPCS_RXCLK_1,
       EPCS_RXDATA,
       EPCS_RXIDLE,
       EPCS_RXRSTN,
       EPCS_RXVAL,
       EPCS_TXCLK,
       EPCS_TXCLK_0,
       EPCS_TXCLK_1,
       EPCS_TXRSTN,
       FATC_RESET_N,
       H2FCALIB0,
       H2FCALIB1,
       M2_ARADDR,
       M2_ARBURST,
       M2_ARID,
       M2_ARLEN,
       M2_ARSIZE,
       M2_ARVALID,
       M2_AWADDR_HADDR,
       M2_AWBURST_HTRANS,
       M2_AWID,
       M2_AWLEN_HBURST,
       M2_AWSIZE_HSIZE,
       M2_AWVALID_HWRITE,
       M2_BREADY,
       M2_RREADY,
       M2_WDATA_HWDATA,
       M2_WID,
       M2_WLAST,
       M2_WSTRB,
       M2_WVALID,
       M_ARADDR,
       M_ARBURST,
       M_ARID,
       M_ARLEN,
       M_ARSIZE,
       M_ARVALID,
       M_AWADDR_HADDR,
       M_AWBURST_HTRANS,
       M_AWID,
       M_AWLEN_HBURST,
       M_AWSIZE_HSIZE,
       M_AWVALID_HWRITE,
       M_BREADY,
       M_RREADY,
       M_WDATA_HWDATA,
       M_WID,
       M_WLAST,
       M_WSTRB,
       M_WVALID,
       PCIE2_LTSSM,
       PCIE2_SYSTEM_INT,
       PCIE2_WAKE_N,
       PCIE_LTSSM,
       PCIE_SYSTEM_INT,
       PLL_LOCK_INT,
       PLL_LOCKLOST_INT,
       S2_ARREADY,
       S2_AWREADY,
       S2_BID,
       S2_BRESP_HRESP,
       S2_BVALID,
       S2_RDATA_HRDATA,
       S2_RID,
       S2_RLAST,
       S2_RRESP,
       S2_RVALID,
       S2_WREADY_HREADYOUT,
       S_ARREADY,
       S_AWREADY,
       S_BID,
       S_BRESP_HRESP,
       S_BVALID,
       S_RDATA_HRDATA,
       S_RID,
       S_RLAST,
       S_RRESP,
       S_RVALID,
       S_WREADY_HREADYOUT,
       SPLL_LOCK,
       WAKE_N,
       XAUI_OUT_CLK,
       APB_CLK,
       APB_PADDR,
       APB_PENABLE,
       APB_PSEL,
       APB_PWDATA,
       APB_PWRITE,
       APB_RSTN,
       CLK_BASE,
       EPCS_PWRDN,
       EPCS_RSTN,
       EPCS_RXERR,
       EPCS_TXDATA,
       EPCS_TXOOB,
       EPCS_TXVAL,
       F2HCALIB0,
       F2HCALIB1,
       FAB_PLL_LOCK,
       FAB_REF_CLK,
       M2_ARREADY,
       M2_AWREADY,
       M2_BID,
       M2_BRESP_HRESP,
       M2_BVALID,
       M2_RDATA_HRDATA,
       M2_RID,
       M2_RLAST,
       M2_RRESP,
       M2_RVALID,
       M2_WREADY_HREADY,
       M_ARREADY,
       M_AWREADY,
       M_BID,
       M_BRESP_HRESP,
       M_BVALID,
       M_RDATA_HRDATA,
       M_RID,
       M_RLAST,
       M_RRESP,
       M_RVALID,
       M_WREADY_HREADY,
       PCIE2_INTERRUPT,
       PCIE2_PERST_N,
       PCIE2_SERDESIF_CORE_RESET_N,
       PCIE2_WAKE_REQ,
       PCIE_INTERRUPT,
       PERST_N,
       S2_ARADDR,
       S2_ARBURST,
       S2_ARID,
       S2_ARLEN,
       S2_ARLOCK,
       S2_ARSIZE,
       S2_ARVALID,
       S2_AWADDR_HADDR,
       S2_AWBURST_HTRANS,
       S2_AWID_HSEL,
       S2_AWLEN_HBURST,
       S2_AWLOCK,
       S2_AWSIZE_HSIZE,
       S2_AWVALID_HWRITE,
       S2_BREADY_HREADY,
       S2_RREADY,
       S2_WDATA_HWDATA,
       S2_WID,
       S2_WLAST,
       S2_WSTRB,
       S2_WVALID,
       S_ARADDR,
       S_ARBURST,
       S_ARID,
       S_ARLEN,
       S_ARLOCK,
       S_ARSIZE,
       S_ARVALID,
       S_AWADDR_HADDR,
       S_AWBURST_HTRANS,
       S_AWID_HSEL,
       S_AWLEN_HBURST,
       S_AWLOCK,
       S_AWSIZE_HSIZE,
       S_AWVALID_HWRITE,
       S_BREADY_HREADY,
       S_RREADY,
       S_WDATA_HWDATA,
       S_WID,
       S_WLAST,
       S_WSTRB,
       S_WVALID,
       SERDESIF_CORE_RESET_N,
       SERDESIF_PHY_RESET_N,
       WAKE_REQ,
       XAUI_FB_CLK,
       RXD3_P,
       RXD2_P,
       RXD1_P,
       RXD0_P,
       RXD3_N,
       RXD2_N,
       RXD1_N,
       RXD0_N,
       TXD3_P,
       TXD2_P,
       TXD1_P,
       TXD0_P,
       TXD3_N,
       TXD2_N,
       TXD1_N,
       TXD0_N,
       REFCLK0,
       REFCLK1
    ) ;
/* synthesis syn_black_box

syn_tsu0 = " APB_PADDR[10]->APB_CLK = 3.791"
syn_tsu1 = " APB_PADDR[11]->APB_CLK = 3.498"
syn_tsu2 = " APB_PADDR[12]->APB_CLK = 3.309"
syn_tsu3 = " APB_PADDR[13]->APB_CLK = 3.076"
syn_tsu4 = " APB_PADDR[14]->APB_CLK = 2.521"
syn_tsu5 = " APB_PADDR[2]->APB_CLK = 2.929"
syn_tsu6 = " APB_PADDR[3]->APB_CLK = 3.244"
syn_tsu7 = " APB_PADDR[4]->APB_CLK = 2.893"
syn_tsu8 = " APB_PADDR[5]->APB_CLK = 3.29"
syn_tsu9 = " APB_PADDR[6]->APB_CLK = 2.853"
syn_tsu10 = " APB_PADDR[7]->APB_CLK = 2.851"
syn_tsu11 = " APB_PADDR[8]->APB_CLK = 3.48"
syn_tsu12 = " APB_PADDR[9]->APB_CLK = 3.473"
syn_tsu13 = " APB_PENABLE->APB_CLK = 0.833"
syn_tsu14 = " APB_PSEL->APB_CLK = 2.83"
syn_tsu15 = " APB_PWDATA[0]->APB_CLK = 1.294"
syn_tsu16 = " APB_PWDATA[10]->APB_CLK = 0.494"
syn_tsu17 = " APB_PWDATA[11]->APB_CLK = 0.581"
syn_tsu18 = " APB_PWDATA[12]->APB_CLK = 0.831"
syn_tsu19 = " APB_PWDATA[13]->APB_CLK = 0.725"
syn_tsu20 = " APB_PWDATA[14]->APB_CLK = 0.897"
syn_tsu21 = " APB_PWDATA[15]->APB_CLK = 0.713"
syn_tsu22 = " APB_PWDATA[16]->APB_CLK = 0.813"
syn_tsu23 = " APB_PWDATA[17]->APB_CLK = 0.747"
syn_tsu24 = " APB_PWDATA[18]->APB_CLK = 0.748"
syn_tsu25 = " APB_PWDATA[19]->APB_CLK = 0.954"
syn_tsu26 = " APB_PWDATA[1]->APB_CLK = 1.879"
syn_tsu27 = " APB_PWDATA[20]->APB_CLK = 0.803"
syn_tsu28 = " APB_PWDATA[21]->APB_CLK = 0.46"
syn_tsu29 = " APB_PWDATA[22]->APB_CLK = 0.516"
syn_tsu30 = " APB_PWDATA[23]->APB_CLK = 0.496"
syn_tsu31 = " APB_PWDATA[24]->APB_CLK = 0.642"
syn_tsu32 = " APB_PWDATA[25]->APB_CLK = 0.509"
syn_tsu33 = " APB_PWDATA[26]->APB_CLK = 0.421"
syn_tsu34 = " APB_PWDATA[27]->APB_CLK = 0.546"
syn_tsu35 = " APB_PWDATA[28]->APB_CLK = 0.087"
syn_tsu36 = " APB_PWDATA[29]->APB_CLK = 0"
syn_tsu37 = " APB_PWDATA[2]->APB_CLK = 1.743"
syn_tsu38 = " APB_PWDATA[30]->APB_CLK = 0.556"
syn_tsu39 = " APB_PWDATA[31]->APB_CLK = 0.054"
syn_tsu40 = " APB_PWDATA[3]->APB_CLK = 1.95"
syn_tsu41 = " APB_PWDATA[4]->APB_CLK = 1.925"
syn_tsu42 = " APB_PWDATA[5]->APB_CLK = 1.226"
syn_tsu43 = " APB_PWDATA[6]->APB_CLK = 1.954"
syn_tsu44 = " APB_PWDATA[7]->APB_CLK = 0.928"
syn_tsu45 = " APB_PWDATA[8]->APB_CLK = 0.693"
syn_tsu46 = " APB_PWDATA[9]->APB_CLK = 0.849"
syn_tsu47 = " APB_PWRITE->APB_CLK = 1.751"
syn_tsu48 = " M2_ARREADY->CLK_BASE = 0.92"
syn_tsu49 = " M2_AWREADY->CLK_BASE = 0.812"
syn_tsu50 = " M2_BID[0]->CLK_BASE = 0.079"
syn_tsu51 = " M2_BRESP_HRESP[0]->CLK_BASE = 0.119"
syn_tsu52 = " M2_BVALID->CLK_BASE = 0.892"
syn_tsu53 = " M2_RDATA_HRDATA[0]->CLK_BASE = 0.632"
syn_tsu54 = " M2_RDATA_HRDATA[10]->CLK_BASE = 0.666"
syn_tsu55 = " M2_RDATA_HRDATA[11]->CLK_BASE = 0.53"
syn_tsu56 = " M2_RDATA_HRDATA[12]->CLK_BASE = 0.706"
syn_tsu57 = " M2_RDATA_HRDATA[13]->CLK_BASE = 0.283"
syn_tsu58 = " M2_RDATA_HRDATA[14]->CLK_BASE = 0.626"
syn_tsu59 = " M2_RDATA_HRDATA[15]->CLK_BASE = 0.499"
syn_tsu60 = " M2_RDATA_HRDATA[16]->CLK_BASE = 0.761"
syn_tsu61 = " M2_RDATA_HRDATA[17]->CLK_BASE = 0.529"
syn_tsu62 = " M2_RDATA_HRDATA[18]->CLK_BASE = 0.721"
syn_tsu63 = " M2_RDATA_HRDATA[19]->CLK_BASE = 0.751"
syn_tsu64 = " M2_RDATA_HRDATA[1]->CLK_BASE = 0.691"
syn_tsu65 = " M2_RDATA_HRDATA[20]->CLK_BASE = 0.417"
syn_tsu66 = " M2_RDATA_HRDATA[21]->CLK_BASE = 0.449"
syn_tsu67 = " M2_RDATA_HRDATA[22]->CLK_BASE = 0.28"
syn_tsu68 = " M2_RDATA_HRDATA[23]->CLK_BASE = 0.657"
syn_tsu69 = " M2_RDATA_HRDATA[24]->CLK_BASE = 0.75"
syn_tsu70 = " M2_RDATA_HRDATA[25]->CLK_BASE = 0.841"
syn_tsu71 = " M2_RDATA_HRDATA[26]->CLK_BASE = 0.572"
syn_tsu72 = " M2_RDATA_HRDATA[27]->CLK_BASE = 0.174"
syn_tsu73 = " M2_RDATA_HRDATA[28]->CLK_BASE = 0.712"
syn_tsu74 = " M2_RDATA_HRDATA[29]->CLK_BASE = 0.707"
syn_tsu75 = " M2_RDATA_HRDATA[2]->CLK_BASE = 0.769"
syn_tsu76 = " M2_RDATA_HRDATA[30]->CLK_BASE = 0.389"
syn_tsu77 = " M2_RDATA_HRDATA[31]->CLK_BASE = 0.729"
syn_tsu78 = " M2_RDATA_HRDATA[32]->CLK_BASE = 0.879"
syn_tsu79 = " M2_RDATA_HRDATA[33]->CLK_BASE = 0.853"
syn_tsu80 = " M2_RDATA_HRDATA[34]->CLK_BASE = 0"
syn_tsu81 = " M2_RDATA_HRDATA[35]->CLK_BASE = 0.191"
syn_tsu82 = " M2_RDATA_HRDATA[36]->CLK_BASE = 0.532"
syn_tsu83 = " M2_RDATA_HRDATA[37]->CLK_BASE = 0.525"
syn_tsu84 = " M2_RDATA_HRDATA[38]->CLK_BASE = 0.953"
syn_tsu85 = " M2_RDATA_HRDATA[39]->CLK_BASE = 0.458"
syn_tsu86 = " M2_RDATA_HRDATA[3]->CLK_BASE = 0.83"
syn_tsu87 = " M2_RDATA_HRDATA[40]->CLK_BASE = 0.557"
syn_tsu88 = " M2_RDATA_HRDATA[41]->CLK_BASE = 0.571"
syn_tsu89 = " M2_RDATA_HRDATA[42]->CLK_BASE = 0.379"
syn_tsu90 = " M2_RDATA_HRDATA[43]->CLK_BASE = 0.795"
syn_tsu91 = " M2_RDATA_HRDATA[44]->CLK_BASE = 0.942"
syn_tsu92 = " M2_RDATA_HRDATA[45]->CLK_BASE = 0.537"
syn_tsu93 = " M2_RDATA_HRDATA[46]->CLK_BASE = 0.791"
syn_tsu94 = " M2_RDATA_HRDATA[47]->CLK_BASE = 0.021"
syn_tsu95 = " M2_RDATA_HRDATA[48]->CLK_BASE = 0.436"
syn_tsu96 = " M2_RDATA_HRDATA[49]->CLK_BASE = 0.803"
syn_tsu97 = " M2_RDATA_HRDATA[4]->CLK_BASE = 0.53"
syn_tsu98 = " M2_RDATA_HRDATA[50]->CLK_BASE = 0.186"
syn_tsu99 = " M2_RDATA_HRDATA[51]->CLK_BASE = 0.894"
syn_tsu100 = " M2_RDATA_HRDATA[52]->CLK_BASE = 0.495"
syn_tsu101 = " M2_RDATA_HRDATA[53]->CLK_BASE = 0.649"
syn_tsu102 = " M2_RDATA_HRDATA[54]->CLK_BASE = 0.518"
syn_tsu103 = " M2_RDATA_HRDATA[55]->CLK_BASE = 0.62"
syn_tsu104 = " M2_RDATA_HRDATA[56]->CLK_BASE = 0.717"
syn_tsu105 = " M2_RDATA_HRDATA[57]->CLK_BASE = 0.69"
syn_tsu106 = " M2_RDATA_HRDATA[58]->CLK_BASE = 0.589"
syn_tsu107 = " M2_RDATA_HRDATA[59]->CLK_BASE = 0.927"
syn_tsu108 = " M2_RDATA_HRDATA[5]->CLK_BASE = 0.58"
syn_tsu109 = " M2_RDATA_HRDATA[60]->CLK_BASE = 0.524"
syn_tsu110 = " M2_RDATA_HRDATA[61]->CLK_BASE = 0.329"
syn_tsu111 = " M2_RDATA_HRDATA[62]->CLK_BASE = 0.598"
syn_tsu112 = " M2_RDATA_HRDATA[63]->CLK_BASE = 0.822"
syn_tsu113 = " M2_RDATA_HRDATA[6]->CLK_BASE = 0.806"
syn_tsu114 = " M2_RDATA_HRDATA[7]->CLK_BASE = 0.747"
syn_tsu115 = " M2_RDATA_HRDATA[8]->CLK_BASE = 0.325"
syn_tsu116 = " M2_RDATA_HRDATA[9]->CLK_BASE = 0.655"
syn_tsu117 = " M2_RID[0]->CLK_BASE = 0.6"
syn_tsu118 = " M2_RID[1]->CLK_BASE = 0.634"
syn_tsu119 = " M2_RID[2]->CLK_BASE = 0.103"
syn_tsu120 = " M2_RID[3]->CLK_BASE = 0.533"
syn_tsu121 = " M2_RLAST->CLK_BASE = 0.628"
syn_tsu122 = " M2_RRESP[0]->CLK_BASE = 0.216"
syn_tsu123 = " M2_RRESP[1]->CLK_BASE = 0.721"
syn_tsu124 = " M2_RVALID->CLK_BASE = 0.936"
syn_tsu125 = " M2_WREADY_HREADY->CLK_BASE = 0.991"
syn_tsu126 = " M_ARREADY->CLK_BASE = 0.86"
syn_tsu127 = " M_AWREADY->CLK_BASE = 1.008"
syn_tsu128 = " M_BID[0]->CLK_BASE = 0.564"
syn_tsu129 = " M_BRESP_HRESP[0]->CLK_BASE = 0.392"
syn_tsu130 = " M_BVALID->CLK_BASE = 0.596"
syn_tsu131 = " M_RDATA_HRDATA[0]->CLK_BASE = 0.787"
syn_tsu132 = " M_RDATA_HRDATA[10]->CLK_BASE = 0.781"
syn_tsu133 = " M_RDATA_HRDATA[11]->CLK_BASE = 0.977"
syn_tsu134 = " M_RDATA_HRDATA[12]->CLK_BASE = 0.553"
syn_tsu135 = " M_RDATA_HRDATA[13]->CLK_BASE = 0.804"
syn_tsu136 = " M_RDATA_HRDATA[14]->CLK_BASE = 0.605"
syn_tsu137 = " M_RDATA_HRDATA[15]->CLK_BASE = 0.914"
syn_tsu138 = " M_RDATA_HRDATA[16]->CLK_BASE = 0.67"
syn_tsu139 = " M_RDATA_HRDATA[17]->CLK_BASE = 0.579"
syn_tsu140 = " M_RDATA_HRDATA[18]->CLK_BASE = 0.557"
syn_tsu141 = " M_RDATA_HRDATA[19]->CLK_BASE = 0.732"
syn_tsu142 = " M_RDATA_HRDATA[1]->CLK_BASE = 0.748"
syn_tsu143 = " M_RDATA_HRDATA[20]->CLK_BASE = 0.604"
syn_tsu144 = " M_RDATA_HRDATA[21]->CLK_BASE = 0.795"
syn_tsu145 = " M_RDATA_HRDATA[22]->CLK_BASE = 0.96"
syn_tsu146 = " M_RDATA_HRDATA[23]->CLK_BASE = 0.9"
syn_tsu147 = " M_RDATA_HRDATA[24]->CLK_BASE = 0.339"
syn_tsu148 = " M_RDATA_HRDATA[25]->CLK_BASE = 0.755"
syn_tsu149 = " M_RDATA_HRDATA[26]->CLK_BASE = 0.537"
syn_tsu150 = " M_RDATA_HRDATA[27]->CLK_BASE = 0.6"
syn_tsu151 = " M_RDATA_HRDATA[28]->CLK_BASE = 0.771"
syn_tsu152 = " M_RDATA_HRDATA[29]->CLK_BASE = 0.531"
syn_tsu153 = " M_RDATA_HRDATA[2]->CLK_BASE = 0.934"
syn_tsu154 = " M_RDATA_HRDATA[30]->CLK_BASE = 0.567"
syn_tsu155 = " M_RDATA_HRDATA[31]->CLK_BASE = 0.631"
syn_tsu156 = " M_RDATA_HRDATA[32]->CLK_BASE = 0.737"
syn_tsu157 = " M_RDATA_HRDATA[33]->CLK_BASE = 0.538"
syn_tsu158 = " M_RDATA_HRDATA[34]->CLK_BASE = 0.756"
syn_tsu159 = " M_RDATA_HRDATA[35]->CLK_BASE = 0.628"
syn_tsu160 = " M_RDATA_HRDATA[36]->CLK_BASE = 0.282"
syn_tsu161 = " M_RDATA_HRDATA[37]->CLK_BASE = 0.847"
syn_tsu162 = " M_RDATA_HRDATA[38]->CLK_BASE = 0.689"
syn_tsu163 = " M_RDATA_HRDATA[39]->CLK_BASE = 0.941"
syn_tsu164 = " M_RDATA_HRDATA[3]->CLK_BASE = 0.868"
syn_tsu165 = " M_RDATA_HRDATA[40]->CLK_BASE = 0.7"
syn_tsu166 = " M_RDATA_HRDATA[41]->CLK_BASE = 0.798"
syn_tsu167 = " M_RDATA_HRDATA[42]->CLK_BASE = 0.902"
syn_tsu168 = " M_RDATA_HRDATA[43]->CLK_BASE = 0.707"
syn_tsu169 = " M_RDATA_HRDATA[44]->CLK_BASE = 0.877"
syn_tsu170 = " M_RDATA_HRDATA[45]->CLK_BASE = 0.595"
syn_tsu171 = " M_RDATA_HRDATA[46]->CLK_BASE = 0.929"
syn_tsu172 = " M_RDATA_HRDATA[47]->CLK_BASE = 0.827"
syn_tsu173 = " M_RDATA_HRDATA[48]->CLK_BASE = 0.532"
syn_tsu174 = " M_RDATA_HRDATA[49]->CLK_BASE = 0.801"
syn_tsu175 = " M_RDATA_HRDATA[4]->CLK_BASE = 0.734"
syn_tsu176 = " M_RDATA_HRDATA[50]->CLK_BASE = 0.835"
syn_tsu177 = " M_RDATA_HRDATA[51]->CLK_BASE = 0.887"
syn_tsu178 = " M_RDATA_HRDATA[52]->CLK_BASE = 0.889"
syn_tsu179 = " M_RDATA_HRDATA[53]->CLK_BASE = 0.745"
syn_tsu180 = " M_RDATA_HRDATA[54]->CLK_BASE = 0.768"
syn_tsu181 = " M_RDATA_HRDATA[55]->CLK_BASE = 0.607"
syn_tsu182 = " M_RDATA_HRDATA[56]->CLK_BASE = 0.82"
syn_tsu183 = " M_RDATA_HRDATA[57]->CLK_BASE = 0.295"
syn_tsu184 = " M_RDATA_HRDATA[58]->CLK_BASE = 0.414"
syn_tsu185 = " M_RDATA_HRDATA[59]->CLK_BASE = 0.92"
syn_tsu186 = " M_RDATA_HRDATA[5]->CLK_BASE = 0.852"
syn_tsu187 = " M_RDATA_HRDATA[60]->CLK_BASE = 0.448"
syn_tsu188 = " M_RDATA_HRDATA[61]->CLK_BASE = 0.785"
syn_tsu189 = " M_RDATA_HRDATA[62]->CLK_BASE = 0.458"
syn_tsu190 = " M_RDATA_HRDATA[63]->CLK_BASE = 0.884"
syn_tsu191 = " M_RDATA_HRDATA[6]->CLK_BASE = 0.401"
syn_tsu192 = " M_RDATA_HRDATA[7]->CLK_BASE = 0.623"
syn_tsu193 = " M_RDATA_HRDATA[8]->CLK_BASE = 0.911"
syn_tsu194 = " M_RDATA_HRDATA[9]->CLK_BASE = 0.709"
syn_tsu195 = " M_RID[0]->CLK_BASE = 0.596"
syn_tsu196 = " M_RID[1]->CLK_BASE = 0.114"
syn_tsu197 = " M_RID[2]->CLK_BASE = 0.661"
syn_tsu198 = " M_RID[3]->CLK_BASE = 0.561"
syn_tsu199 = " M_RLAST->CLK_BASE = 0.791"
syn_tsu200 = " M_RRESP[0]->CLK_BASE = 0.741"
syn_tsu201 = " M_RRESP[1]->CLK_BASE = 0.53"
syn_tsu202 = " M_RVALID->CLK_BASE = 0.348"
syn_tsu203 = " M_WREADY_HREADY->CLK_BASE = 1.052"
syn_tsu204 = " S2_ARADDR[0]->CLK_BASE = 0.564"
syn_tsu205 = " S2_ARADDR[10]->CLK_BASE = 0.454"
syn_tsu206 = " S2_ARADDR[11]->CLK_BASE = 0.669"
syn_tsu207 = " S2_ARADDR[12]->CLK_BASE = 0.169"
syn_tsu208 = " S2_ARADDR[13]->CLK_BASE = 0.143"
syn_tsu209 = " S2_ARADDR[14]->CLK_BASE = 0.487"
syn_tsu210 = " S2_ARADDR[15]->CLK_BASE = 0.468"
syn_tsu211 = " S2_ARADDR[16]->CLK_BASE = 0.135"
syn_tsu212 = " S2_ARADDR[17]->CLK_BASE = 0.11"
syn_tsu213 = " S2_ARADDR[18]->CLK_BASE = 0.972"
syn_tsu214 = " S2_ARADDR[19]->CLK_BASE = 0.432"
syn_tsu215 = " S2_ARADDR[1]->CLK_BASE = 0.552"
syn_tsu216 = " S2_ARADDR[20]->CLK_BASE = 0.414"
syn_tsu217 = " S2_ARADDR[21]->CLK_BASE = 0.431"
syn_tsu218 = " S2_ARADDR[22]->CLK_BASE = 0.512"
syn_tsu219 = " S2_ARADDR[23]->CLK_BASE = 0.486"
syn_tsu220 = " S2_ARADDR[24]->CLK_BASE = 0.421"
syn_tsu221 = " S2_ARADDR[25]->CLK_BASE = 0.764"
syn_tsu222 = " S2_ARADDR[26]->CLK_BASE = 0.913"
syn_tsu223 = " S2_ARADDR[27]->CLK_BASE = 0.455"
syn_tsu224 = " S2_ARADDR[28]->CLK_BASE = 0.996"
syn_tsu225 = " S2_ARADDR[29]->CLK_BASE = 0.497"
syn_tsu226 = " S2_ARADDR[2]->CLK_BASE = 0.905"
syn_tsu227 = " S2_ARADDR[30]->CLK_BASE = 0.309"
syn_tsu228 = " S2_ARADDR[31]->CLK_BASE = 0.687"
syn_tsu229 = " S2_ARADDR[3]->CLK_BASE = 0.151"
syn_tsu230 = " S2_ARADDR[4]->CLK_BASE = 0.344"
syn_tsu231 = " S2_ARADDR[5]->CLK_BASE = 0.015"
syn_tsu232 = " S2_ARADDR[6]->CLK_BASE = 0.219"
syn_tsu233 = " S2_ARADDR[7]->CLK_BASE = 1.025"
syn_tsu234 = " S2_ARADDR[8]->CLK_BASE = 0.451"
syn_tsu235 = " S2_ARADDR[9]->CLK_BASE = 0.058"
syn_tsu236 = " S2_ARBURST[0]->CLK_BASE = 0.517"
syn_tsu237 = " S2_ARBURST[1]->CLK_BASE = 0.586"
syn_tsu238 = " S2_ARID[0]->CLK_BASE = 0.139"
syn_tsu239 = " S2_ARID[1]->CLK_BASE = 0.243"
syn_tsu240 = " S2_ARID[2]->CLK_BASE = 0.226"
syn_tsu241 = " S2_ARID[3]->CLK_BASE = 0.473"
syn_tsu242 = " S2_ARLEN[0]->CLK_BASE = 0.279"
syn_tsu243 = " S2_ARLEN[1]->CLK_BASE = 0.54"
syn_tsu244 = " S2_ARLEN[2]->CLK_BASE = 0.12"
syn_tsu245 = " S2_ARLEN[3]->CLK_BASE = 0.149"
syn_tsu246 = " S2_ARSIZE[0]->CLK_BASE = 0.885"
syn_tsu247 = " S2_ARSIZE[1]->CLK_BASE = 0.532"
syn_tsu248 = " S2_ARVALID->CLK_BASE = 0.392"
syn_tsu249 = " S2_AWADDR_HADDR[0]->CLK_BASE = 0.721"
syn_tsu250 = " S2_AWADDR_HADDR[10]->CLK_BASE = 0.746"
syn_tsu251 = " S2_AWADDR_HADDR[11]->CLK_BASE = 0.568"
syn_tsu252 = " S2_AWADDR_HADDR[12]->CLK_BASE = 0.257"
syn_tsu253 = " S2_AWADDR_HADDR[13]->CLK_BASE = 0.334"
syn_tsu254 = " S2_AWADDR_HADDR[14]->CLK_BASE = 0.446"
syn_tsu255 = " S2_AWADDR_HADDR[15]->CLK_BASE = 0.294"
syn_tsu256 = " S2_AWADDR_HADDR[16]->CLK_BASE = 0.611"
syn_tsu257 = " S2_AWADDR_HADDR[17]->CLK_BASE = 0.435"
syn_tsu258 = " S2_AWADDR_HADDR[18]->CLK_BASE = 0.843"
syn_tsu259 = " S2_AWADDR_HADDR[19]->CLK_BASE = 0.914"
syn_tsu260 = " S2_AWADDR_HADDR[1]->CLK_BASE = 0.464"
syn_tsu261 = " S2_AWADDR_HADDR[20]->CLK_BASE = 0.448"
syn_tsu262 = " S2_AWADDR_HADDR[21]->CLK_BASE = 0.758"
syn_tsu263 = " S2_AWADDR_HADDR[22]->CLK_BASE = 0.672"
syn_tsu264 = " S2_AWADDR_HADDR[23]->CLK_BASE = 0.845"
syn_tsu265 = " S2_AWADDR_HADDR[24]->CLK_BASE = 0.613"
syn_tsu266 = " S2_AWADDR_HADDR[25]->CLK_BASE = 0.65"
syn_tsu267 = " S2_AWADDR_HADDR[26]->CLK_BASE = 0.75"
syn_tsu268 = " S2_AWADDR_HADDR[27]->CLK_BASE = 0.509"
syn_tsu269 = " S2_AWADDR_HADDR[28]->CLK_BASE = 0.672"
syn_tsu270 = " S2_AWADDR_HADDR[29]->CLK_BASE = 0.409"
syn_tsu271 = " S2_AWADDR_HADDR[2]->CLK_BASE = 0.3"
syn_tsu272 = " S2_AWADDR_HADDR[30]->CLK_BASE = 0.933"
syn_tsu273 = " S2_AWADDR_HADDR[31]->CLK_BASE = 0.87"
syn_tsu274 = " S2_AWADDR_HADDR[3]->CLK_BASE = 0.494"
syn_tsu275 = " S2_AWADDR_HADDR[4]->CLK_BASE = 0.64"
syn_tsu276 = " S2_AWADDR_HADDR[5]->CLK_BASE = 0.326"
syn_tsu277 = " S2_AWADDR_HADDR[6]->CLK_BASE = 0.781"
syn_tsu278 = " S2_AWADDR_HADDR[7]->CLK_BASE = 0.341"
syn_tsu279 = " S2_AWADDR_HADDR[8]->CLK_BASE = 0.838"
syn_tsu280 = " S2_AWADDR_HADDR[9]->CLK_BASE = 0.538"
syn_tsu281 = " S2_AWBURST_HTRANS[0]->CLK_BASE = 0.937"
syn_tsu282 = " S2_AWBURST_HTRANS[1]->CLK_BASE = 1.035"
syn_tsu283 = " S2_AWID_HSEL[0]->CLK_BASE = 1.065"
syn_tsu284 = " S2_AWID_HSEL[1]->CLK_BASE = 0.164"
syn_tsu285 = " S2_AWID_HSEL[2]->CLK_BASE = 0.109"
syn_tsu286 = " S2_AWID_HSEL[3]->CLK_BASE = 0"
syn_tsu287 = " S2_AWLEN_HBURST[0]->CLK_BASE = 0.071"
syn_tsu288 = " S2_AWLEN_HBURST[1]->CLK_BASE = 0"
syn_tsu289 = " S2_AWLEN_HBURST[2]->CLK_BASE = 0.037"
syn_tsu290 = " S2_AWLEN_HBURST[3]->CLK_BASE = 0.425"
syn_tsu291 = " S2_AWSIZE_HSIZE[0]->CLK_BASE = 0.939"
syn_tsu292 = " S2_AWSIZE_HSIZE[1]->CLK_BASE = 0.74"
syn_tsu293 = " S2_AWVALID_HWRITE->CLK_BASE = 0.798"
syn_tsu294 = " S2_BREADY_HREADY->CLK_BASE = 0.972"
syn_tsu295 = " S2_RREADY->CLK_BASE = 0.85"
syn_tsu296 = " S2_WDATA_HWDATA[0]->CLK_BASE = 0.007"
syn_tsu297 = " S2_WDATA_HWDATA[10]->CLK_BASE = 0.147"
syn_tsu298 = " S2_WDATA_HWDATA[11]->CLK_BASE = 0.088"
syn_tsu299 = " S2_WDATA_HWDATA[12]->CLK_BASE = 0.187"
syn_tsu300 = " S2_WDATA_HWDATA[13]->CLK_BASE = 0.242"
syn_tsu301 = " S2_WDATA_HWDATA[14]->CLK_BASE = 0.179"
syn_tsu302 = " S2_WDATA_HWDATA[15]->CLK_BASE = 0.12"
syn_tsu303 = " S2_WDATA_HWDATA[16]->CLK_BASE = 0.108"
syn_tsu304 = " S2_WDATA_HWDATA[17]->CLK_BASE = 0.173"
syn_tsu305 = " S2_WDATA_HWDATA[18]->CLK_BASE = 0.427"
syn_tsu306 = " S2_WDATA_HWDATA[19]->CLK_BASE = 0.236"
syn_tsu307 = " S2_WDATA_HWDATA[1]->CLK_BASE = 0.051"
syn_tsu308 = " S2_WDATA_HWDATA[20]->CLK_BASE = 0.281"
syn_tsu309 = " S2_WDATA_HWDATA[21]->CLK_BASE = 0"
syn_tsu310 = " S2_WDATA_HWDATA[22]->CLK_BASE = 0.144"
syn_tsu311 = " S2_WDATA_HWDATA[23]->CLK_BASE = 0.163"
syn_tsu312 = " S2_WDATA_HWDATA[24]->CLK_BASE = 0.324"
syn_tsu313 = " S2_WDATA_HWDATA[25]->CLK_BASE = 0.307"
syn_tsu314 = " S2_WDATA_HWDATA[26]->CLK_BASE = 0.169"
syn_tsu315 = " S2_WDATA_HWDATA[27]->CLK_BASE = 0.185"
syn_tsu316 = " S2_WDATA_HWDATA[28]->CLK_BASE = 0.436"
syn_tsu317 = " S2_WDATA_HWDATA[29]->CLK_BASE = 0.353"
syn_tsu318 = " S2_WDATA_HWDATA[2]->CLK_BASE = 0.136"
syn_tsu319 = " S2_WDATA_HWDATA[30]->CLK_BASE = 0.152"
syn_tsu320 = " S2_WDATA_HWDATA[31]->CLK_BASE = 0.288"
syn_tsu321 = " S2_WDATA_HWDATA[32]->CLK_BASE = 0.19"
syn_tsu322 = " S2_WDATA_HWDATA[33]->CLK_BASE = 0.555"
syn_tsu323 = " S2_WDATA_HWDATA[34]->CLK_BASE = 0.466"
syn_tsu324 = " S2_WDATA_HWDATA[35]->CLK_BASE = 0.424"
syn_tsu325 = " S2_WDATA_HWDATA[36]->CLK_BASE = 0.212"
syn_tsu326 = " S2_WDATA_HWDATA[37]->CLK_BASE = 0.026"
syn_tsu327 = " S2_WDATA_HWDATA[38]->CLK_BASE = 0.004"
syn_tsu328 = " S2_WDATA_HWDATA[39]->CLK_BASE = 0"
syn_tsu329 = " S2_WDATA_HWDATA[3]->CLK_BASE = 0.044"
syn_tsu330 = " S2_WDATA_HWDATA[40]->CLK_BASE = 0"
syn_tsu331 = " S2_WDATA_HWDATA[41]->CLK_BASE = 0"
syn_tsu332 = " S2_WDATA_HWDATA[42]->CLK_BASE = 0.447"
syn_tsu333 = " S2_WDATA_HWDATA[43]->CLK_BASE = 0.703"
syn_tsu334 = " S2_WDATA_HWDATA[44]->CLK_BASE = 0"
syn_tsu335 = " S2_WDATA_HWDATA[45]->CLK_BASE = 0.037"
syn_tsu336 = " S2_WDATA_HWDATA[46]->CLK_BASE = 0.295"
syn_tsu337 = " S2_WDATA_HWDATA[47]->CLK_BASE = 0"
syn_tsu338 = " S2_WDATA_HWDATA[48]->CLK_BASE = 0.505"
syn_tsu339 = " S2_WDATA_HWDATA[49]->CLK_BASE = 0.176"
syn_tsu340 = " S2_WDATA_HWDATA[4]->CLK_BASE = 0.38"
syn_tsu341 = " S2_WDATA_HWDATA[50]->CLK_BASE = 0.269"
syn_tsu342 = " S2_WDATA_HWDATA[51]->CLK_BASE = 0.11"
syn_tsu343 = " S2_WDATA_HWDATA[52]->CLK_BASE = 0.046"
syn_tsu344 = " S2_WDATA_HWDATA[53]->CLK_BASE = 0"
syn_tsu345 = " S2_WDATA_HWDATA[54]->CLK_BASE = 0.045"
syn_tsu346 = " S2_WDATA_HWDATA[55]->CLK_BASE = 0"
syn_tsu347 = " S2_WDATA_HWDATA[56]->CLK_BASE = 0.423"
syn_tsu348 = " S2_WDATA_HWDATA[57]->CLK_BASE = 0.37"
syn_tsu349 = " S2_WDATA_HWDATA[58]->CLK_BASE = 0.004"
syn_tsu350 = " S2_WDATA_HWDATA[59]->CLK_BASE = 0"
syn_tsu351 = " S2_WDATA_HWDATA[5]->CLK_BASE = 0.432"
syn_tsu352 = " S2_WDATA_HWDATA[60]->CLK_BASE = 0.046"
syn_tsu353 = " S2_WDATA_HWDATA[61]->CLK_BASE = 0"
syn_tsu354 = " S2_WDATA_HWDATA[62]->CLK_BASE = 0.428"
syn_tsu355 = " S2_WDATA_HWDATA[63]->CLK_BASE = 0.148"
syn_tsu356 = " S2_WDATA_HWDATA[6]->CLK_BASE = 0.137"
syn_tsu357 = " S2_WDATA_HWDATA[7]->CLK_BASE = 0.407"
syn_tsu358 = " S2_WDATA_HWDATA[8]->CLK_BASE = 0.669"
syn_tsu359 = " S2_WDATA_HWDATA[9]->CLK_BASE = 0.093"
syn_tsu360 = " S2_WLAST->CLK_BASE = 0.265"
syn_tsu361 = " S2_WSTRB[0]->CLK_BASE = 0.685"
syn_tsu362 = " S2_WSTRB[1]->CLK_BASE = 0.313"
syn_tsu363 = " S2_WSTRB[2]->CLK_BASE = 0.535"
syn_tsu364 = " S2_WSTRB[3]->CLK_BASE = 0.323"
syn_tsu365 = " S2_WSTRB[4]->CLK_BASE = 0.083"
syn_tsu366 = " S2_WSTRB[5]->CLK_BASE = 0.671"
syn_tsu367 = " S2_WSTRB[6]->CLK_BASE = 0.424"
syn_tsu368 = " S2_WSTRB[7]->CLK_BASE = 0.391"
syn_tsu369 = " S2_WVALID->CLK_BASE = 0.437"
syn_tsu370 = " S_ARADDR[0]->CLK_BASE = 0.852"
syn_tsu371 = " S_ARADDR[10]->CLK_BASE = 1.011"
syn_tsu372 = " S_ARADDR[11]->CLK_BASE = 0.989"
syn_tsu373 = " S_ARADDR[12]->CLK_BASE = 0.622"
syn_tsu374 = " S_ARADDR[13]->CLK_BASE = 0.694"
syn_tsu375 = " S_ARADDR[14]->CLK_BASE = 0.938"
syn_tsu376 = " S_ARADDR[15]->CLK_BASE = 0.545"
syn_tsu377 = " S_ARADDR[16]->CLK_BASE = 0.513"
syn_tsu378 = " S_ARADDR[17]->CLK_BASE = 0.871"
syn_tsu379 = " S_ARADDR[18]->CLK_BASE = 1.032"
syn_tsu380 = " S_ARADDR[19]->CLK_BASE = 0.883"
syn_tsu381 = " S_ARADDR[1]->CLK_BASE = 0.42"
syn_tsu382 = " S_ARADDR[20]->CLK_BASE = 0.873"
syn_tsu383 = " S_ARADDR[21]->CLK_BASE = 0.757"
syn_tsu384 = " S_ARADDR[22]->CLK_BASE = 0.761"
syn_tsu385 = " S_ARADDR[23]->CLK_BASE = 0.942"
syn_tsu386 = " S_ARADDR[24]->CLK_BASE = 0.556"
syn_tsu387 = " S_ARADDR[25]->CLK_BASE = 0.594"
syn_tsu388 = " S_ARADDR[26]->CLK_BASE = 0.599"
syn_tsu389 = " S_ARADDR[27]->CLK_BASE = 0.923"
syn_tsu390 = " S_ARADDR[28]->CLK_BASE = 0.588"
syn_tsu391 = " S_ARADDR[29]->CLK_BASE = 0.713"
syn_tsu392 = " S_ARADDR[2]->CLK_BASE = 0.736"
syn_tsu393 = " S_ARADDR[30]->CLK_BASE = 0.68"
syn_tsu394 = " S_ARADDR[31]->CLK_BASE = 0.659"
syn_tsu395 = " S_ARADDR[3]->CLK_BASE = 1.077"
syn_tsu396 = " S_ARADDR[4]->CLK_BASE = 0.514"
syn_tsu397 = " S_ARADDR[5]->CLK_BASE = 0.678"
syn_tsu398 = " S_ARADDR[6]->CLK_BASE = 1.054"
syn_tsu399 = " S_ARADDR[7]->CLK_BASE = 0.686"
syn_tsu400 = " S_ARADDR[8]->CLK_BASE = 0.971"
syn_tsu401 = " S_ARADDR[9]->CLK_BASE = 0.791"
syn_tsu402 = " S_ARBURST[0]->CLK_BASE = 0.564"
syn_tsu403 = " S_ARBURST[1]->CLK_BASE = 0.491"
syn_tsu404 = " S_ARID[0]->CLK_BASE = 0.656"
syn_tsu405 = " S_ARID[1]->CLK_BASE = 0.647"
syn_tsu406 = " S_ARID[2]->CLK_BASE = 0.708"
syn_tsu407 = " S_ARID[3]->CLK_BASE = 0.638"
syn_tsu408 = " S_ARLEN[0]->CLK_BASE = 0.569"
syn_tsu409 = " S_ARLEN[1]->CLK_BASE = 0.659"
syn_tsu410 = " S_ARLEN[2]->CLK_BASE = 0.607"
syn_tsu411 = " S_ARLEN[3]->CLK_BASE = 0.511"
syn_tsu412 = " S_ARSIZE[0]->CLK_BASE = 0.618"
syn_tsu413 = " S_ARSIZE[1]->CLK_BASE = 0.896"
syn_tsu414 = " S_ARVALID->CLK_BASE = 0.664"
syn_tsu415 = " S_AWADDR_HADDR[0]->CLK_BASE = 0.622"
syn_tsu416 = " S_AWADDR_HADDR[10]->CLK_BASE = 0.797"
syn_tsu417 = " S_AWADDR_HADDR[11]->CLK_BASE = 0.933"
syn_tsu418 = " S_AWADDR_HADDR[12]->CLK_BASE = 0.739"
syn_tsu419 = " S_AWADDR_HADDR[13]->CLK_BASE = 0.878"
syn_tsu420 = " S_AWADDR_HADDR[14]->CLK_BASE = 0.821"
syn_tsu421 = " S_AWADDR_HADDR[15]->CLK_BASE = 0.614"
syn_tsu422 = " S_AWADDR_HADDR[16]->CLK_BASE = 0.704"
syn_tsu423 = " S_AWADDR_HADDR[17]->CLK_BASE = 0.839"
syn_tsu424 = " S_AWADDR_HADDR[18]->CLK_BASE = 1.037"
syn_tsu425 = " S_AWADDR_HADDR[19]->CLK_BASE = 0.748"
syn_tsu426 = " S_AWADDR_HADDR[1]->CLK_BASE = 0.677"
syn_tsu427 = " S_AWADDR_HADDR[20]->CLK_BASE = 0.727"
syn_tsu428 = " S_AWADDR_HADDR[21]->CLK_BASE = 0.819"
syn_tsu429 = " S_AWADDR_HADDR[22]->CLK_BASE = 0.886"
syn_tsu430 = " S_AWADDR_HADDR[23]->CLK_BASE = 0.76"
syn_tsu431 = " S_AWADDR_HADDR[24]->CLK_BASE = 0.63"
syn_tsu432 = " S_AWADDR_HADDR[25]->CLK_BASE = 0.972"
syn_tsu433 = " S_AWADDR_HADDR[26]->CLK_BASE = 0.513"
syn_tsu434 = " S_AWADDR_HADDR[27]->CLK_BASE = 0.89"
syn_tsu435 = " S_AWADDR_HADDR[28]->CLK_BASE = 0.67"
syn_tsu436 = " S_AWADDR_HADDR[29]->CLK_BASE = 0.9"
syn_tsu437 = " S_AWADDR_HADDR[2]->CLK_BASE = 0.612"
syn_tsu438 = " S_AWADDR_HADDR[30]->CLK_BASE = 0.884"
syn_tsu439 = " S_AWADDR_HADDR[31]->CLK_BASE = 0.751"
syn_tsu440 = " S_AWADDR_HADDR[3]->CLK_BASE = 0.924"
syn_tsu441 = " S_AWADDR_HADDR[4]->CLK_BASE = 0.584"
syn_tsu442 = " S_AWADDR_HADDR[5]->CLK_BASE = 0.479"
syn_tsu443 = " S_AWADDR_HADDR[6]->CLK_BASE = 0.65"
syn_tsu444 = " S_AWADDR_HADDR[7]->CLK_BASE = 0.937"
syn_tsu445 = " S_AWADDR_HADDR[8]->CLK_BASE = 0.454"
syn_tsu446 = " S_AWADDR_HADDR[9]->CLK_BASE = 0.665"
syn_tsu447 = " S_AWBURST_HTRANS[0]->CLK_BASE = 0.862"
syn_tsu448 = " S_AWBURST_HTRANS[1]->CLK_BASE = 0.881"
syn_tsu449 = " S_AWID_HSEL[0]->CLK_BASE = 0.793"
syn_tsu450 = " S_AWID_HSEL[1]->CLK_BASE = 0.46"
syn_tsu451 = " S_AWID_HSEL[2]->CLK_BASE = 0.422"
syn_tsu452 = " S_AWID_HSEL[3]->CLK_BASE = 0.245"
syn_tsu453 = " S_AWLEN_HBURST[0]->CLK_BASE = 0.53"
syn_tsu454 = " S_AWLEN_HBURST[1]->CLK_BASE = 0.207"
syn_tsu455 = " S_AWLEN_HBURST[2]->CLK_BASE = 0.582"
syn_tsu456 = " S_AWLEN_HBURST[3]->CLK_BASE = 0.649"
syn_tsu457 = " S_AWSIZE_HSIZE[0]->CLK_BASE = 0.996"
syn_tsu458 = " S_AWSIZE_HSIZE[1]->CLK_BASE = 0.963"
syn_tsu459 = " S_AWVALID_HWRITE->CLK_BASE = 0.783"
syn_tsu460 = " S_BREADY_HREADY->CLK_BASE = 1.046"
syn_tsu461 = " S_RREADY->CLK_BASE = 0.878"
syn_tsu462 = " S_WDATA_HWDATA[0]->CLK_BASE = 0.548"
syn_tsu463 = " S_WDATA_HWDATA[10]->CLK_BASE = 0.273"
syn_tsu464 = " S_WDATA_HWDATA[11]->CLK_BASE = 0.544"
syn_tsu465 = " S_WDATA_HWDATA[12]->CLK_BASE = 0.351"
syn_tsu466 = " S_WDATA_HWDATA[13]->CLK_BASE = 0.607"
syn_tsu467 = " S_WDATA_HWDATA[14]->CLK_BASE = 0.284"
syn_tsu468 = " S_WDATA_HWDATA[15]->CLK_BASE = 0.328"
syn_tsu469 = " S_WDATA_HWDATA[16]->CLK_BASE = 0.379"
syn_tsu470 = " S_WDATA_HWDATA[17]->CLK_BASE = 0.668"
syn_tsu471 = " S_WDATA_HWDATA[18]->CLK_BASE = 0.496"
syn_tsu472 = " S_WDATA_HWDATA[19]->CLK_BASE = 0.333"
syn_tsu473 = " S_WDATA_HWDATA[1]->CLK_BASE = 0.646"
syn_tsu474 = " S_WDATA_HWDATA[20]->CLK_BASE = 0.381"
syn_tsu475 = " S_WDATA_HWDATA[21]->CLK_BASE = 0.462"
syn_tsu476 = " S_WDATA_HWDATA[22]->CLK_BASE = 0.32"
syn_tsu477 = " S_WDATA_HWDATA[23]->CLK_BASE = 0.621"
syn_tsu478 = " S_WDATA_HWDATA[24]->CLK_BASE = 0.258"
syn_tsu479 = " S_WDATA_HWDATA[25]->CLK_BASE = 0.38"
syn_tsu480 = " S_WDATA_HWDATA[26]->CLK_BASE = 0.529"
syn_tsu481 = " S_WDATA_HWDATA[27]->CLK_BASE = 0.659"
syn_tsu482 = " S_WDATA_HWDATA[28]->CLK_BASE = 0.334"
syn_tsu483 = " S_WDATA_HWDATA[29]->CLK_BASE = 0.546"
syn_tsu484 = " S_WDATA_HWDATA[2]->CLK_BASE = 0.241"
syn_tsu485 = " S_WDATA_HWDATA[30]->CLK_BASE = 0.245"
syn_tsu486 = " S_WDATA_HWDATA[31]->CLK_BASE = 0.684"
syn_tsu487 = " S_WDATA_HWDATA[32]->CLK_BASE = 0.658"
syn_tsu488 = " S_WDATA_HWDATA[33]->CLK_BASE = 0.712"
syn_tsu489 = " S_WDATA_HWDATA[34]->CLK_BASE = 0.726"
syn_tsu490 = " S_WDATA_HWDATA[35]->CLK_BASE = 0.756"
syn_tsu491 = " S_WDATA_HWDATA[36]->CLK_BASE = 0.301"
syn_tsu492 = " S_WDATA_HWDATA[37]->CLK_BASE = 0.562"
syn_tsu493 = " S_WDATA_HWDATA[38]->CLK_BASE = 0.715"
syn_tsu494 = " S_WDATA_HWDATA[39]->CLK_BASE = 0.52"
syn_tsu495 = " S_WDATA_HWDATA[3]->CLK_BASE = 0.288"
syn_tsu496 = " S_WDATA_HWDATA[40]->CLK_BASE = 0.297"
syn_tsu497 = " S_WDATA_HWDATA[41]->CLK_BASE = 0.524"
syn_tsu498 = " S_WDATA_HWDATA[42]->CLK_BASE = 0.723"
syn_tsu499 = " S_WDATA_HWDATA[43]->CLK_BASE = 0.715"
syn_tsu500 = " S_WDATA_HWDATA[44]->CLK_BASE = 0.353"
syn_tsu501 = " S_WDATA_HWDATA[45]->CLK_BASE = 0.349"
syn_tsu502 = " S_WDATA_HWDATA[46]->CLK_BASE = 0.783"
syn_tsu503 = " S_WDATA_HWDATA[47]->CLK_BASE = 0.467"
syn_tsu504 = " S_WDATA_HWDATA[48]->CLK_BASE = 0.519"
syn_tsu505 = " S_WDATA_HWDATA[49]->CLK_BASE = 0.336"
syn_tsu506 = " S_WDATA_HWDATA[4]->CLK_BASE = 0.231"
syn_tsu507 = " S_WDATA_HWDATA[50]->CLK_BASE = 0.34"
syn_tsu508 = " S_WDATA_HWDATA[51]->CLK_BASE = 0.747"
syn_tsu509 = " S_WDATA_HWDATA[52]->CLK_BASE = 0.578"
syn_tsu510 = " S_WDATA_HWDATA[53]->CLK_BASE = 0.664"
syn_tsu511 = " S_WDATA_HWDATA[54]->CLK_BASE = 0.69"
syn_tsu512 = " S_WDATA_HWDATA[55]->CLK_BASE = 0.567"
syn_tsu513 = " S_WDATA_HWDATA[56]->CLK_BASE = 0.752"
syn_tsu514 = " S_WDATA_HWDATA[57]->CLK_BASE = 0.56"
syn_tsu515 = " S_WDATA_HWDATA[58]->CLK_BASE = 0.541"
syn_tsu516 = " S_WDATA_HWDATA[59]->CLK_BASE = 0.487"
syn_tsu517 = " S_WDATA_HWDATA[5]->CLK_BASE = 0.253"
syn_tsu518 = " S_WDATA_HWDATA[60]->CLK_BASE = 0.58"
syn_tsu519 = " S_WDATA_HWDATA[61]->CLK_BASE = 0.552"
syn_tsu520 = " S_WDATA_HWDATA[62]->CLK_BASE = 0.291"
syn_tsu521 = " S_WDATA_HWDATA[63]->CLK_BASE = 0.53"
syn_tsu522 = " S_WDATA_HWDATA[6]->CLK_BASE = 0.631"
syn_tsu523 = " S_WDATA_HWDATA[7]->CLK_BASE = 0.726"
syn_tsu524 = " S_WDATA_HWDATA[8]->CLK_BASE = 0.303"
syn_tsu525 = " S_WDATA_HWDATA[9]->CLK_BASE = 0.32"
syn_tsu526 = " S_WLAST->CLK_BASE = 0.467"
syn_tsu527 = " S_WSTRB[0]->CLK_BASE = 0.711"
syn_tsu528 = " S_WSTRB[1]->CLK_BASE = 0.827"
syn_tsu529 = " S_WSTRB[2]->CLK_BASE = 0.955"
syn_tsu530 = " S_WSTRB[3]->CLK_BASE = 0.862"
syn_tsu531 = " S_WSTRB[4]->CLK_BASE = 0.537"
syn_tsu532 = " S_WSTRB[5]->CLK_BASE = 0.91"
syn_tsu533 = " S_WSTRB[6]->CLK_BASE = 0.403"
syn_tsu534 = " S_WSTRB[7]->CLK_BASE = 0.633"
syn_tsu535 = " S_WVALID->CLK_BASE = 0.703"
syn_tco0 = " APB_CLK->APB_PRDATA[0] = 4.934"
syn_tco1 = " APB_CLK->APB_PRDATA[10] = 5.024"
syn_tco2 = " APB_CLK->APB_PRDATA[11] = 5.105"
syn_tco3 = " APB_CLK->APB_PRDATA[12] = 5.156"
syn_tco4 = " APB_CLK->APB_PRDATA[13] = 5.196"
syn_tco5 = " APB_CLK->APB_PRDATA[14] = 5.014"
syn_tco6 = " APB_CLK->APB_PRDATA[15] = 5.106"
syn_tco7 = " APB_CLK->APB_PRDATA[16] = 5.048"
syn_tco8 = " APB_CLK->APB_PRDATA[17] = 5.201"
syn_tco9 = " APB_CLK->APB_PRDATA[18] = 5.007"
syn_tco10 = " APB_CLK->APB_PRDATA[19] = 5.160"
syn_tco11 = " APB_CLK->APB_PRDATA[1] = 4.896"
syn_tco12 = " APB_CLK->APB_PRDATA[20] = 5.049"
syn_tco13 = " APB_CLK->APB_PRDATA[21] = 5.157"
syn_tco14 = " APB_CLK->APB_PRDATA[22] = 5.029"
syn_tco15 = " APB_CLK->APB_PRDATA[23] = 5.161"
syn_tco16 = " APB_CLK->APB_PRDATA[24] = 5.230"
syn_tco17 = " APB_CLK->APB_PRDATA[25] = 5.348"
syn_tco18 = " APB_CLK->APB_PRDATA[26] = 5.076"
syn_tco19 = " APB_CLK->APB_PRDATA[27] = 5.125"
syn_tco20 = " APB_CLK->APB_PRDATA[28] = 5.217"
syn_tco21 = " APB_CLK->APB_PRDATA[29] = 5.235"
syn_tco22 = " APB_CLK->APB_PRDATA[2] = 5.014"
syn_tco23 = " APB_CLK->APB_PRDATA[30] = 4.986"
syn_tco24 = " APB_CLK->APB_PRDATA[31] = 5.038"
syn_tco25 = " APB_CLK->APB_PRDATA[3] = 4.838"
syn_tco26 = " APB_CLK->APB_PRDATA[4] = 4.918"
syn_tco27 = " APB_CLK->APB_PRDATA[5] = 4.908"
syn_tco28 = " APB_CLK->APB_PRDATA[6] = 4.814"
syn_tco29 = " APB_CLK->APB_PRDATA[7] = 4.869"
syn_tco30 = " APB_CLK->APB_PRDATA[8] = 5.255"
syn_tco31 = " APB_CLK->APB_PRDATA[9] = 5.129"
syn_tco32 = " APB_CLK->APB_PREADY = 4.732"
syn_tco33 = " APB_CLK->APB_PSLVERR = 4.957"
syn_tco34 = " APB_CLK->PCIE2_SYSTEM_INT = 3.792"
syn_tco35 = " APB_CLK->PCIE_SYSTEM_INT = 4.040"
syn_tco36 = " APB_CLK->PLL_LOCKLOST_INT = 3.655"
syn_tco37 = " APB_CLK->PLL_LOCK_INT = 3.873"
syn_tco38 = " CLK_BASE->M2_ARADDR[0] = 3.154"
syn_tco39 = " CLK_BASE->M2_ARADDR[10] = 3.207"
syn_tco40 = " CLK_BASE->M2_ARADDR[11] = 3.120"
syn_tco41 = " CLK_BASE->M2_ARADDR[12] = 3.218"
syn_tco42 = " CLK_BASE->M2_ARADDR[13] = 3.227"
syn_tco43 = " CLK_BASE->M2_ARADDR[14] = 3.268"
syn_tco44 = " CLK_BASE->M2_ARADDR[15] = 3.253"
syn_tco45 = " CLK_BASE->M2_ARADDR[16] = 3.215"
syn_tco46 = " CLK_BASE->M2_ARADDR[17] = 3.229"
syn_tco47 = " CLK_BASE->M2_ARADDR[18] = 3.184"
syn_tco48 = " CLK_BASE->M2_ARADDR[19] = 3.181"
syn_tco49 = " CLK_BASE->M2_ARADDR[1] = 3.133"
syn_tco50 = " CLK_BASE->M2_ARADDR[20] = 3.125"
syn_tco51 = " CLK_BASE->M2_ARADDR[21] = 3.251"
syn_tco52 = " CLK_BASE->M2_ARADDR[22] = 3.190"
syn_tco53 = " CLK_BASE->M2_ARADDR[23] = 3.229"
syn_tco54 = " CLK_BASE->M2_ARADDR[24] = 3.238"
syn_tco55 = " CLK_BASE->M2_ARADDR[25] = 3.071"
syn_tco56 = " CLK_BASE->M2_ARADDR[26] = 3.105"
syn_tco57 = " CLK_BASE->M2_ARADDR[27] = 3.206"
syn_tco58 = " CLK_BASE->M2_ARADDR[28] = 3.191"
syn_tco59 = " CLK_BASE->M2_ARADDR[29] = 3.127"
syn_tco60 = " CLK_BASE->M2_ARADDR[2] = 3.180"
syn_tco61 = " CLK_BASE->M2_ARADDR[30] = 3.080"
syn_tco62 = " CLK_BASE->M2_ARADDR[31] = 3.207"
syn_tco63 = " CLK_BASE->M2_ARADDR[3] = 3.130"
syn_tco64 = " CLK_BASE->M2_ARADDR[4] = 3.135"
syn_tco65 = " CLK_BASE->M2_ARADDR[5] = 3.116"
syn_tco66 = " CLK_BASE->M2_ARADDR[6] = 3.218"
syn_tco67 = " CLK_BASE->M2_ARADDR[7] = 3.150"
syn_tco68 = " CLK_BASE->M2_ARADDR[8] = 3.163"
syn_tco69 = " CLK_BASE->M2_ARADDR[9] = 3.256"
syn_tco70 = " CLK_BASE->M2_ARBURST[0] = 3.128"
syn_tco71 = " CLK_BASE->M2_ARID[0] = 3.117"
syn_tco72 = " CLK_BASE->M2_ARID[1] = 3.094"
syn_tco73 = " CLK_BASE->M2_ARLEN[0] = 3.156"
syn_tco74 = " CLK_BASE->M2_ARLEN[1] = 3.137"
syn_tco75 = " CLK_BASE->M2_ARLEN[2] = 3.086"
syn_tco76 = " CLK_BASE->M2_ARLEN[3] = 3.112"
syn_tco77 = " CLK_BASE->M2_ARSIZE[0] = 3.176"
syn_tco78 = " CLK_BASE->M2_ARSIZE[1] = 3.161"
syn_tco79 = " CLK_BASE->M2_ARVALID = 3.171"
syn_tco80 = " CLK_BASE->M2_AWADDR_HADDR[10] = 3.057"
syn_tco81 = " CLK_BASE->M2_AWADDR_HADDR[11] = 3.038"
syn_tco82 = " CLK_BASE->M2_AWADDR_HADDR[12] = 3.093"
syn_tco83 = " CLK_BASE->M2_AWADDR_HADDR[13] = 3.040"
syn_tco84 = " CLK_BASE->M2_AWADDR_HADDR[14] = 3.051"
syn_tco85 = " CLK_BASE->M2_AWADDR_HADDR[15] = 3.105"
syn_tco86 = " CLK_BASE->M2_AWADDR_HADDR[16] = 3.087"
syn_tco87 = " CLK_BASE->M2_AWADDR_HADDR[17] = 3.095"
syn_tco88 = " CLK_BASE->M2_AWADDR_HADDR[18] = 3.123"
syn_tco89 = " CLK_BASE->M2_AWADDR_HADDR[19] = 3.057"
syn_tco90 = " CLK_BASE->M2_AWADDR_HADDR[20] = 3.167"
syn_tco91 = " CLK_BASE->M2_AWADDR_HADDR[21] = 3.124"
syn_tco92 = " CLK_BASE->M2_AWADDR_HADDR[22] = 3.054"
syn_tco93 = " CLK_BASE->M2_AWADDR_HADDR[23] = 3.033"
syn_tco94 = " CLK_BASE->M2_AWADDR_HADDR[24] = 3.125"
syn_tco95 = " CLK_BASE->M2_AWADDR_HADDR[25] = 3.047"
syn_tco96 = " CLK_BASE->M2_AWADDR_HADDR[26] = 3.076"
syn_tco97 = " CLK_BASE->M2_AWADDR_HADDR[27] = 3.046"
syn_tco98 = " CLK_BASE->M2_AWADDR_HADDR[28] = 3.058"
syn_tco99 = " CLK_BASE->M2_AWADDR_HADDR[29] = 3.215"
syn_tco100 = " CLK_BASE->M2_AWADDR_HADDR[2] = 3.132"
syn_tco101 = " CLK_BASE->M2_AWADDR_HADDR[30] = 3.168"
syn_tco102 = " CLK_BASE->M2_AWADDR_HADDR[31] = 3.035"
syn_tco103 = " CLK_BASE->M2_AWADDR_HADDR[3] = 3.181"
syn_tco104 = " CLK_BASE->M2_AWADDR_HADDR[4] = 3.044"
syn_tco105 = " CLK_BASE->M2_AWADDR_HADDR[5] = 3.242"
syn_tco106 = " CLK_BASE->M2_AWADDR_HADDR[6] = 3.248"
syn_tco107 = " CLK_BASE->M2_AWADDR_HADDR[7] = 3.182"
syn_tco108 = " CLK_BASE->M2_AWADDR_HADDR[8] = 3.239"
syn_tco109 = " CLK_BASE->M2_AWADDR_HADDR[9] = 3.035"
syn_tco110 = " CLK_BASE->M2_AWBURST_HTRANS[0] = 3.188"
syn_tco111 = " CLK_BASE->M2_AWLEN_HBURST[0] = 3.007"
syn_tco112 = " CLK_BASE->M2_AWLEN_HBURST[1] = 3.010"
syn_tco113 = " CLK_BASE->M2_AWLEN_HBURST[2] = 3.006"
syn_tco114 = " CLK_BASE->M2_AWLEN_HBURST[3] = 3.035"
syn_tco115 = " CLK_BASE->M2_AWSIZE_HSIZE[0] = 3.064"
syn_tco116 = " CLK_BASE->M2_AWSIZE_HSIZE[1] = 3.026"
syn_tco117 = " CLK_BASE->M2_AWVALID_HWRITE = 3.190"
syn_tco118 = " CLK_BASE->M2_BREADY = 3.185"
syn_tco119 = " CLK_BASE->M2_RREADY = 2.845"
syn_tco120 = " CLK_BASE->M2_WDATA_HWDATA[0] = 3.172"
syn_tco121 = " CLK_BASE->M2_WDATA_HWDATA[10] = 3.234"
syn_tco122 = " CLK_BASE->M2_WDATA_HWDATA[11] = 3.271"
syn_tco123 = " CLK_BASE->M2_WDATA_HWDATA[12] = 3.269"
syn_tco124 = " CLK_BASE->M2_WDATA_HWDATA[13] = 3.185"
syn_tco125 = " CLK_BASE->M2_WDATA_HWDATA[14] = 3.244"
syn_tco126 = " CLK_BASE->M2_WDATA_HWDATA[15] = 3.234"
syn_tco127 = " CLK_BASE->M2_WDATA_HWDATA[16] = 3.248"
syn_tco128 = " CLK_BASE->M2_WDATA_HWDATA[17] = 3.137"
syn_tco129 = " CLK_BASE->M2_WDATA_HWDATA[18] = 3.193"
syn_tco130 = " CLK_BASE->M2_WDATA_HWDATA[19] = 3.145"
syn_tco131 = " CLK_BASE->M2_WDATA_HWDATA[1] = 3.150"
syn_tco132 = " CLK_BASE->M2_WDATA_HWDATA[20] = 3.141"
syn_tco133 = " CLK_BASE->M2_WDATA_HWDATA[21] = 3.190"
syn_tco134 = " CLK_BASE->M2_WDATA_HWDATA[22] = 3.111"
syn_tco135 = " CLK_BASE->M2_WDATA_HWDATA[23] = 3.109"
syn_tco136 = " CLK_BASE->M2_WDATA_HWDATA[24] = 3.156"
syn_tco137 = " CLK_BASE->M2_WDATA_HWDATA[25] = 3.176"
syn_tco138 = " CLK_BASE->M2_WDATA_HWDATA[26] = 3.153"
syn_tco139 = " CLK_BASE->M2_WDATA_HWDATA[27] = 3.146"
syn_tco140 = " CLK_BASE->M2_WDATA_HWDATA[28] = 3.146"
syn_tco141 = " CLK_BASE->M2_WDATA_HWDATA[29] = 3.250"
syn_tco142 = " CLK_BASE->M2_WDATA_HWDATA[2] = 3.152"
syn_tco143 = " CLK_BASE->M2_WDATA_HWDATA[30] = 3.199"
syn_tco144 = " CLK_BASE->M2_WDATA_HWDATA[31] = 3.120"
syn_tco145 = " CLK_BASE->M2_WDATA_HWDATA[32] = 3.163"
syn_tco146 = " CLK_BASE->M2_WDATA_HWDATA[33] = 3.155"
syn_tco147 = " CLK_BASE->M2_WDATA_HWDATA[34] = 3.148"
syn_tco148 = " CLK_BASE->M2_WDATA_HWDATA[35] = 3.191"
syn_tco149 = " CLK_BASE->M2_WDATA_HWDATA[36] = 3.093"
syn_tco150 = " CLK_BASE->M2_WDATA_HWDATA[37] = 3.198"
syn_tco151 = " CLK_BASE->M2_WDATA_HWDATA[38] = 3.195"
syn_tco152 = " CLK_BASE->M2_WDATA_HWDATA[39] = 3.183"
syn_tco153 = " CLK_BASE->M2_WDATA_HWDATA[3] = 3.197"
syn_tco154 = " CLK_BASE->M2_WDATA_HWDATA[40] = 3.230"
syn_tco155 = " CLK_BASE->M2_WDATA_HWDATA[41] = 3.093"
syn_tco156 = " CLK_BASE->M2_WDATA_HWDATA[42] = 3.165"
syn_tco157 = " CLK_BASE->M2_WDATA_HWDATA[43] = 3.219"
syn_tco158 = " CLK_BASE->M2_WDATA_HWDATA[44] = 3.148"
syn_tco159 = " CLK_BASE->M2_WDATA_HWDATA[45] = 3.183"
syn_tco160 = " CLK_BASE->M2_WDATA_HWDATA[46] = 3.234"
syn_tco161 = " CLK_BASE->M2_WDATA_HWDATA[47] = 3.108"
syn_tco162 = " CLK_BASE->M2_WDATA_HWDATA[48] = 3.255"
syn_tco163 = " CLK_BASE->M2_WDATA_HWDATA[49] = 3.150"
syn_tco164 = " CLK_BASE->M2_WDATA_HWDATA[4] = 3.168"
syn_tco165 = " CLK_BASE->M2_WDATA_HWDATA[50] = 3.163"
syn_tco166 = " CLK_BASE->M2_WDATA_HWDATA[51] = 3.097"
syn_tco167 = " CLK_BASE->M2_WDATA_HWDATA[52] = 3.070"
syn_tco168 = " CLK_BASE->M2_WDATA_HWDATA[53] = 3.190"
syn_tco169 = " CLK_BASE->M2_WDATA_HWDATA[54] = 3.206"
syn_tco170 = " CLK_BASE->M2_WDATA_HWDATA[55] = 3.117"
syn_tco171 = " CLK_BASE->M2_WDATA_HWDATA[56] = 3.193"
syn_tco172 = " CLK_BASE->M2_WDATA_HWDATA[57] = 3.102"
syn_tco173 = " CLK_BASE->M2_WDATA_HWDATA[58] = 3.073"
syn_tco174 = " CLK_BASE->M2_WDATA_HWDATA[59] = 3.082"
syn_tco175 = " CLK_BASE->M2_WDATA_HWDATA[5] = 3.139"
syn_tco176 = " CLK_BASE->M2_WDATA_HWDATA[60] = 3.185"
syn_tco177 = " CLK_BASE->M2_WDATA_HWDATA[61] = 3.144"
syn_tco178 = " CLK_BASE->M2_WDATA_HWDATA[62] = 3.190"
syn_tco179 = " CLK_BASE->M2_WDATA_HWDATA[63] = 3.145"
syn_tco180 = " CLK_BASE->M2_WDATA_HWDATA[6] = 3.214"
syn_tco181 = " CLK_BASE->M2_WDATA_HWDATA[7] = 3.172"
syn_tco182 = " CLK_BASE->M2_WDATA_HWDATA[8] = 3.170"
syn_tco183 = " CLK_BASE->M2_WDATA_HWDATA[9] = 3.104"
syn_tco184 = " CLK_BASE->M2_WLAST = 3.097"
syn_tco185 = " CLK_BASE->M2_WSTRB[0] = 3.174"
syn_tco186 = " CLK_BASE->M2_WSTRB[1] = 3.168"
syn_tco187 = " CLK_BASE->M2_WSTRB[2] = 3.249"
syn_tco188 = " CLK_BASE->M2_WSTRB[3] = 3.145"
syn_tco189 = " CLK_BASE->M2_WSTRB[4] = 3.294"
syn_tco190 = " CLK_BASE->M2_WSTRB[5] = 3.129"
syn_tco191 = " CLK_BASE->M2_WSTRB[6] = 3.172"
syn_tco192 = " CLK_BASE->M2_WSTRB[7] = 3.080"
syn_tco193 = " CLK_BASE->M2_WVALID = 3.207"
syn_tco194 = " CLK_BASE->M_ARADDR[0] = 3.191"
syn_tco195 = " CLK_BASE->M_ARADDR[10] = 3.072"
syn_tco196 = " CLK_BASE->M_ARADDR[11] = 3.066"
syn_tco197 = " CLK_BASE->M_ARADDR[12] = 3.025"
syn_tco198 = " CLK_BASE->M_ARADDR[13] = 3.099"
syn_tco199 = " CLK_BASE->M_ARADDR[14] = 3.006"
syn_tco200 = " CLK_BASE->M_ARADDR[15] = 3.037"
syn_tco201 = " CLK_BASE->M_ARADDR[16] = 3.112"
syn_tco202 = " CLK_BASE->M_ARADDR[17] = 3.007"
syn_tco203 = " CLK_BASE->M_ARADDR[18] = 3.168"
syn_tco204 = " CLK_BASE->M_ARADDR[19] = 3.079"
syn_tco205 = " CLK_BASE->M_ARADDR[1] = 3.211"
syn_tco206 = " CLK_BASE->M_ARADDR[20] = 3.197"
syn_tco207 = " CLK_BASE->M_ARADDR[21] = 3.144"
syn_tco208 = " CLK_BASE->M_ARADDR[22] = 3.163"
syn_tco209 = " CLK_BASE->M_ARADDR[23] = 3.196"
syn_tco210 = " CLK_BASE->M_ARADDR[24] = 3.074"
syn_tco211 = " CLK_BASE->M_ARADDR[25] = 3.147"
syn_tco212 = " CLK_BASE->M_ARADDR[26] = 3.006"
syn_tco213 = " CLK_BASE->M_ARADDR[27] = 2.989"
syn_tco214 = " CLK_BASE->M_ARADDR[28] = 3.130"
syn_tco215 = " CLK_BASE->M_ARADDR[29] = 3.033"
syn_tco216 = " CLK_BASE->M_ARADDR[2] = 3.204"
syn_tco217 = " CLK_BASE->M_ARADDR[30] = 3.071"
syn_tco218 = " CLK_BASE->M_ARADDR[31] = 3.175"
syn_tco219 = " CLK_BASE->M_ARADDR[3] = 3.195"
syn_tco220 = " CLK_BASE->M_ARADDR[4] = 3.021"
syn_tco221 = " CLK_BASE->M_ARADDR[5] = 3.038"
syn_tco222 = " CLK_BASE->M_ARADDR[6] = 3.003"
syn_tco223 = " CLK_BASE->M_ARADDR[7] = 3.061"
syn_tco224 = " CLK_BASE->M_ARADDR[8] = 2.969"
syn_tco225 = " CLK_BASE->M_ARADDR[9] = 3.015"
syn_tco226 = " CLK_BASE->M_ARBURST[0] = 2.990"
syn_tco227 = " CLK_BASE->M_ARID[0] = 2.933"
syn_tco228 = " CLK_BASE->M_ARID[1] = 3.165"
syn_tco229 = " CLK_BASE->M_ARLEN[0] = 2.909"
syn_tco230 = " CLK_BASE->M_ARLEN[1] = 3.087"
syn_tco231 = " CLK_BASE->M_ARLEN[2] = 3.050"
syn_tco232 = " CLK_BASE->M_ARLEN[3] = 2.966"
syn_tco233 = " CLK_BASE->M_ARSIZE[0] = 3.154"
syn_tco234 = " CLK_BASE->M_ARSIZE[1] = 3.170"
syn_tco235 = " CLK_BASE->M_ARVALID = 3.163"
syn_tco236 = " CLK_BASE->M_AWADDR_HADDR[10] = 3.118"
syn_tco237 = " CLK_BASE->M_AWADDR_HADDR[11] = 3.061"
syn_tco238 = " CLK_BASE->M_AWADDR_HADDR[12] = 2.992"
syn_tco239 = " CLK_BASE->M_AWADDR_HADDR[13] = 3.002"
syn_tco240 = " CLK_BASE->M_AWADDR_HADDR[14] = 3.046"
syn_tco241 = " CLK_BASE->M_AWADDR_HADDR[15] = 2.916"
syn_tco242 = " CLK_BASE->M_AWADDR_HADDR[16] = 3.030"
syn_tco243 = " CLK_BASE->M_AWADDR_HADDR[17] = 2.982"
syn_tco244 = " CLK_BASE->M_AWADDR_HADDR[18] = 3.009"
syn_tco245 = " CLK_BASE->M_AWADDR_HADDR[19] = 3.051"
syn_tco246 = " CLK_BASE->M_AWADDR_HADDR[20] = 3.011"
syn_tco247 = " CLK_BASE->M_AWADDR_HADDR[21] = 3.062"
syn_tco248 = " CLK_BASE->M_AWADDR_HADDR[22] = 2.973"
syn_tco249 = " CLK_BASE->M_AWADDR_HADDR[23] = 3.059"
syn_tco250 = " CLK_BASE->M_AWADDR_HADDR[24] = 3.049"
syn_tco251 = " CLK_BASE->M_AWADDR_HADDR[25] = 2.884"
syn_tco252 = " CLK_BASE->M_AWADDR_HADDR[26] = 2.839"
syn_tco253 = " CLK_BASE->M_AWADDR_HADDR[27] = 3.070"
syn_tco254 = " CLK_BASE->M_AWADDR_HADDR[28] = 2.827"
syn_tco255 = " CLK_BASE->M_AWADDR_HADDR[29] = 3.016"
syn_tco256 = " CLK_BASE->M_AWADDR_HADDR[2] = 3.090"
syn_tco257 = " CLK_BASE->M_AWADDR_HADDR[30] = 2.824"
syn_tco258 = " CLK_BASE->M_AWADDR_HADDR[31] = 3.068"
syn_tco259 = " CLK_BASE->M_AWADDR_HADDR[3] = 3.139"
syn_tco260 = " CLK_BASE->M_AWADDR_HADDR[4] = 2.902"
syn_tco261 = " CLK_BASE->M_AWADDR_HADDR[5] = 2.863"
syn_tco262 = " CLK_BASE->M_AWADDR_HADDR[6] = 3.000"
syn_tco263 = " CLK_BASE->M_AWADDR_HADDR[7] = 3.103"
syn_tco264 = " CLK_BASE->M_AWADDR_HADDR[8] = 2.932"
syn_tco265 = " CLK_BASE->M_AWADDR_HADDR[9] = 3.033"
syn_tco266 = " CLK_BASE->M_AWBURST_HTRANS[0] = 2.946"
syn_tco267 = " CLK_BASE->M_AWLEN_HBURST[0] = 3.046"
syn_tco268 = " CLK_BASE->M_AWLEN_HBURST[1] = 3.008"
syn_tco269 = " CLK_BASE->M_AWLEN_HBURST[2] = 2.848"
syn_tco270 = " CLK_BASE->M_AWLEN_HBURST[3] = 2.964"
syn_tco271 = " CLK_BASE->M_AWSIZE_HSIZE[0] = 3.026"
syn_tco272 = " CLK_BASE->M_AWSIZE_HSIZE[1] = 2.902"
syn_tco273 = " CLK_BASE->M_AWVALID_HWRITE = 3.046"
syn_tco274 = " CLK_BASE->M_BREADY = 2.742"
syn_tco275 = " CLK_BASE->M_RREADY = 3.100"
syn_tco276 = " CLK_BASE->M_WDATA_HWDATA[0] = 3.746"
syn_tco277 = " CLK_BASE->M_WDATA_HWDATA[10] = 4.000"
syn_tco278 = " CLK_BASE->M_WDATA_HWDATA[11] = 3.531"
syn_tco279 = " CLK_BASE->M_WDATA_HWDATA[12] = 3.870"
syn_tco280 = " CLK_BASE->M_WDATA_HWDATA[13] = 3.741"
syn_tco281 = " CLK_BASE->M_WDATA_HWDATA[14] = 3.770"
syn_tco282 = " CLK_BASE->M_WDATA_HWDATA[15] = 3.868"
syn_tco283 = " CLK_BASE->M_WDATA_HWDATA[16] = 3.822"
syn_tco284 = " CLK_BASE->M_WDATA_HWDATA[17] = 3.808"
syn_tco285 = " CLK_BASE->M_WDATA_HWDATA[18] = 3.574"
syn_tco286 = " CLK_BASE->M_WDATA_HWDATA[19] = 3.982"
syn_tco287 = " CLK_BASE->M_WDATA_HWDATA[1] = 3.500"
syn_tco288 = " CLK_BASE->M_WDATA_HWDATA[20] = 3.893"
syn_tco289 = " CLK_BASE->M_WDATA_HWDATA[21] = 3.755"
syn_tco290 = " CLK_BASE->M_WDATA_HWDATA[22] = 3.780"
syn_tco291 = " CLK_BASE->M_WDATA_HWDATA[23] = 3.517"
syn_tco292 = " CLK_BASE->M_WDATA_HWDATA[24] = 3.710"
syn_tco293 = " CLK_BASE->M_WDATA_HWDATA[25] = 3.607"
syn_tco294 = " CLK_BASE->M_WDATA_HWDATA[26] = 3.583"
syn_tco295 = " CLK_BASE->M_WDATA_HWDATA[27] = 3.540"
syn_tco296 = " CLK_BASE->M_WDATA_HWDATA[28] = 3.547"
syn_tco297 = " CLK_BASE->M_WDATA_HWDATA[29] = 3.697"
syn_tco298 = " CLK_BASE->M_WDATA_HWDATA[2] = 3.859"
syn_tco299 = " CLK_BASE->M_WDATA_HWDATA[30] = 3.528"
syn_tco300 = " CLK_BASE->M_WDATA_HWDATA[31] = 3.316"
syn_tco301 = " CLK_BASE->M_WDATA_HWDATA[32] = 3.433"
syn_tco302 = " CLK_BASE->M_WDATA_HWDATA[33] = 3.408"
syn_tco303 = " CLK_BASE->M_WDATA_HWDATA[34] = 3.210"
syn_tco304 = " CLK_BASE->M_WDATA_HWDATA[35] = 3.448"
syn_tco305 = " CLK_BASE->M_WDATA_HWDATA[36] = 3.297"
syn_tco306 = " CLK_BASE->M_WDATA_HWDATA[37] = 3.214"
syn_tco307 = " CLK_BASE->M_WDATA_HWDATA[38] = 3.290"
syn_tco308 = " CLK_BASE->M_WDATA_HWDATA[39] = 3.256"
syn_tco309 = " CLK_BASE->M_WDATA_HWDATA[3] = 3.869"
syn_tco310 = " CLK_BASE->M_WDATA_HWDATA[40] = 3.252"
syn_tco311 = " CLK_BASE->M_WDATA_HWDATA[41] = 3.362"
syn_tco312 = " CLK_BASE->M_WDATA_HWDATA[42] = 3.435"
syn_tco313 = " CLK_BASE->M_WDATA_HWDATA[43] = 3.448"
syn_tco314 = " CLK_BASE->M_WDATA_HWDATA[44] = 3.283"
syn_tco315 = " CLK_BASE->M_WDATA_HWDATA[45] = 3.458"
syn_tco316 = " CLK_BASE->M_WDATA_HWDATA[46] = 3.312"
syn_tco317 = " CLK_BASE->M_WDATA_HWDATA[47] = 3.530"
syn_tco318 = " CLK_BASE->M_WDATA_HWDATA[48] = 3.379"
syn_tco319 = " CLK_BASE->M_WDATA_HWDATA[49] = 3.323"
syn_tco320 = " CLK_BASE->M_WDATA_HWDATA[4] = 3.846"
syn_tco321 = " CLK_BASE->M_WDATA_HWDATA[50] = 3.320"
syn_tco322 = " CLK_BASE->M_WDATA_HWDATA[51] = 3.452"
syn_tco323 = " CLK_BASE->M_WDATA_HWDATA[52] = 3.666"
syn_tco324 = " CLK_BASE->M_WDATA_HWDATA[53] = 3.846"
syn_tco325 = " CLK_BASE->M_WDATA_HWDATA[54] = 3.682"
syn_tco326 = " CLK_BASE->M_WDATA_HWDATA[55] = 3.489"
syn_tco327 = " CLK_BASE->M_WDATA_HWDATA[56] = 3.628"
syn_tco328 = " CLK_BASE->M_WDATA_HWDATA[57] = 3.583"
syn_tco329 = " CLK_BASE->M_WDATA_HWDATA[58] = 3.502"
syn_tco330 = " CLK_BASE->M_WDATA_HWDATA[59] = 3.729"
syn_tco331 = " CLK_BASE->M_WDATA_HWDATA[5] = 3.708"
syn_tco332 = " CLK_BASE->M_WDATA_HWDATA[60] = 3.535"
syn_tco333 = " CLK_BASE->M_WDATA_HWDATA[61] = 3.626"
syn_tco334 = " CLK_BASE->M_WDATA_HWDATA[62] = 3.781"
syn_tco335 = " CLK_BASE->M_WDATA_HWDATA[63] = 3.621"
syn_tco336 = " CLK_BASE->M_WDATA_HWDATA[6] = 3.684"
syn_tco337 = " CLK_BASE->M_WDATA_HWDATA[7] = 3.796"
syn_tco338 = " CLK_BASE->M_WDATA_HWDATA[8] = 3.568"
syn_tco339 = " CLK_BASE->M_WDATA_HWDATA[9] = 3.651"
syn_tco340 = " CLK_BASE->M_WLAST = 3.108"
syn_tco341 = " CLK_BASE->M_WSTRB[0] = 3.237"
syn_tco342 = " CLK_BASE->M_WSTRB[1] = 3.676"
syn_tco343 = " CLK_BASE->M_WSTRB[2] = 3.572"
syn_tco344 = " CLK_BASE->M_WSTRB[3] = 3.481"
syn_tco345 = " CLK_BASE->M_WSTRB[4] = 3.574"
syn_tco346 = " CLK_BASE->M_WSTRB[5] = 3.608"
syn_tco347 = " CLK_BASE->M_WSTRB[6] = 3.429"
syn_tco348 = " CLK_BASE->M_WSTRB[7] = 3.575"
syn_tco349 = " CLK_BASE->M_WVALID = 3.090"
syn_tco350 = " CLK_BASE->S2_ARREADY = 3.099"
syn_tco351 = " CLK_BASE->S2_AWREADY = 3.067"
syn_tco352 = " CLK_BASE->S2_BID[0] = 3.109"
syn_tco353 = " CLK_BASE->S2_BID[1] = 3.104"
syn_tco354 = " CLK_BASE->S2_BID[2] = 3.086"
syn_tco355 = " CLK_BASE->S2_BID[3] = 3.045"
syn_tco356 = " CLK_BASE->S2_BRESP_HRESP[1] = 3.194"
syn_tco357 = " CLK_BASE->S2_BVALID = 3.152"
syn_tco358 = " CLK_BASE->S2_RDATA_HRDATA[0] = 3.001"
syn_tco359 = " CLK_BASE->S2_RDATA_HRDATA[10] = 3.047"
syn_tco360 = " CLK_BASE->S2_RDATA_HRDATA[11] = 3.066"
syn_tco361 = " CLK_BASE->S2_RDATA_HRDATA[12] = 3.070"
syn_tco362 = " CLK_BASE->S2_RDATA_HRDATA[13] = 3.017"
syn_tco363 = " CLK_BASE->S2_RDATA_HRDATA[14] = 3.034"
syn_tco364 = " CLK_BASE->S2_RDATA_HRDATA[15] = 3.016"
syn_tco365 = " CLK_BASE->S2_RDATA_HRDATA[16] = 3.039"
syn_tco366 = " CLK_BASE->S2_RDATA_HRDATA[17] = 3.015"
syn_tco367 = " CLK_BASE->S2_RDATA_HRDATA[18] = 3.000"
syn_tco368 = " CLK_BASE->S2_RDATA_HRDATA[19] = 3.023"
syn_tco369 = " CLK_BASE->S2_RDATA_HRDATA[1] = 2.991"
syn_tco370 = " CLK_BASE->S2_RDATA_HRDATA[20] = 3.045"
syn_tco371 = " CLK_BASE->S2_RDATA_HRDATA[21] = 3.006"
syn_tco372 = " CLK_BASE->S2_RDATA_HRDATA[22] = 3.019"
syn_tco373 = " CLK_BASE->S2_RDATA_HRDATA[23] = 3.014"
syn_tco374 = " CLK_BASE->S2_RDATA_HRDATA[24] = 3.018"
syn_tco375 = " CLK_BASE->S2_RDATA_HRDATA[25] = 3.058"
syn_tco376 = " CLK_BASE->S2_RDATA_HRDATA[26] = 3.003"
syn_tco377 = " CLK_BASE->S2_RDATA_HRDATA[27] = 3.108"
syn_tco378 = " CLK_BASE->S2_RDATA_HRDATA[28] = 3.010"
syn_tco379 = " CLK_BASE->S2_RDATA_HRDATA[29] = 2.980"
syn_tco380 = " CLK_BASE->S2_RDATA_HRDATA[2] = 2.986"
syn_tco381 = " CLK_BASE->S2_RDATA_HRDATA[30] = 2.964"
syn_tco382 = " CLK_BASE->S2_RDATA_HRDATA[31] = 3.098"
syn_tco383 = " CLK_BASE->S2_RDATA_HRDATA[32] = 3.044"
syn_tco384 = " CLK_BASE->S2_RDATA_HRDATA[33] = 3.175"
syn_tco385 = " CLK_BASE->S2_RDATA_HRDATA[34] = 3.131"
syn_tco386 = " CLK_BASE->S2_RDATA_HRDATA[35] = 3.105"
syn_tco387 = " CLK_BASE->S2_RDATA_HRDATA[36] = 3.146"
syn_tco388 = " CLK_BASE->S2_RDATA_HRDATA[37] = 3.101"
syn_tco389 = " CLK_BASE->S2_RDATA_HRDATA[38] = 3.026"
syn_tco390 = " CLK_BASE->S2_RDATA_HRDATA[39] = 3.134"
syn_tco391 = " CLK_BASE->S2_RDATA_HRDATA[3] = 2.967"
syn_tco392 = " CLK_BASE->S2_RDATA_HRDATA[40] = 3.147"
syn_tco393 = " CLK_BASE->S2_RDATA_HRDATA[41] = 3.089"
syn_tco394 = " CLK_BASE->S2_RDATA_HRDATA[42] = 3.145"
syn_tco395 = " CLK_BASE->S2_RDATA_HRDATA[43] = 3.139"
syn_tco396 = " CLK_BASE->S2_RDATA_HRDATA[44] = 3.086"
syn_tco397 = " CLK_BASE->S2_RDATA_HRDATA[45] = 3.174"
syn_tco398 = " CLK_BASE->S2_RDATA_HRDATA[46] = 3.178"
syn_tco399 = " CLK_BASE->S2_RDATA_HRDATA[47] = 3.119"
syn_tco400 = " CLK_BASE->S2_RDATA_HRDATA[48] = 3.172"
syn_tco401 = " CLK_BASE->S2_RDATA_HRDATA[49] = 3.060"
syn_tco402 = " CLK_BASE->S2_RDATA_HRDATA[4] = 3.052"
syn_tco403 = " CLK_BASE->S2_RDATA_HRDATA[50] = 3.157"
syn_tco404 = " CLK_BASE->S2_RDATA_HRDATA[51] = 3.117"
syn_tco405 = " CLK_BASE->S2_RDATA_HRDATA[52] = 3.175"
syn_tco406 = " CLK_BASE->S2_RDATA_HRDATA[53] = 3.053"
syn_tco407 = " CLK_BASE->S2_RDATA_HRDATA[54] = 3.111"
syn_tco408 = " CLK_BASE->S2_RDATA_HRDATA[55] = 3.064"
syn_tco409 = " CLK_BASE->S2_RDATA_HRDATA[56] = 3.159"
syn_tco410 = " CLK_BASE->S2_RDATA_HRDATA[57] = 3.093"
syn_tco411 = " CLK_BASE->S2_RDATA_HRDATA[58] = 3.150"
syn_tco412 = " CLK_BASE->S2_RDATA_HRDATA[59] = 3.088"
syn_tco413 = " CLK_BASE->S2_RDATA_HRDATA[5] = 3.082"
syn_tco414 = " CLK_BASE->S2_RDATA_HRDATA[60] = 3.101"
syn_tco415 = " CLK_BASE->S2_RDATA_HRDATA[61] = 3.029"
syn_tco416 = " CLK_BASE->S2_RDATA_HRDATA[62] = 2.968"
syn_tco417 = " CLK_BASE->S2_RDATA_HRDATA[63] = 3.044"
syn_tco418 = " CLK_BASE->S2_RDATA_HRDATA[6] = 3.065"
syn_tco419 = " CLK_BASE->S2_RDATA_HRDATA[7] = 3.012"
syn_tco420 = " CLK_BASE->S2_RDATA_HRDATA[8] = 3.036"
syn_tco421 = " CLK_BASE->S2_RDATA_HRDATA[9] = 3.005"
syn_tco422 = " CLK_BASE->S2_RID[0] = 2.927"
syn_tco423 = " CLK_BASE->S2_RID[1] = 3.011"
syn_tco424 = " CLK_BASE->S2_RID[2] = 3.018"
syn_tco425 = " CLK_BASE->S2_RID[3] = 2.942"
syn_tco426 = " CLK_BASE->S2_RLAST = 3.084"
syn_tco427 = " CLK_BASE->S2_RRESP[1] = 2.948"
syn_tco428 = " CLK_BASE->S2_RVALID = 3.161"
syn_tco429 = " CLK_BASE->S2_WREADY_HREADYOUT = 2.645"
syn_tco430 = " CLK_BASE->S_ARREADY = 2.901"
syn_tco431 = " CLK_BASE->S_AWREADY = 2.934"
syn_tco432 = " CLK_BASE->S_BID[0] = 3.098"
syn_tco433 = " CLK_BASE->S_BID[1] = 3.147"
syn_tco434 = " CLK_BASE->S_BID[2] = 3.169"
syn_tco435 = " CLK_BASE->S_BID[3] = 3.215"
syn_tco436 = " CLK_BASE->S_BRESP_HRESP[1] = 3.199"
syn_tco437 = " CLK_BASE->S_BVALID = 3.251"
syn_tco438 = " CLK_BASE->S_RDATA_HRDATA[0] = 3.170"
syn_tco439 = " CLK_BASE->S_RDATA_HRDATA[10] = 3.148"
syn_tco440 = " CLK_BASE->S_RDATA_HRDATA[11] = 3.170"
syn_tco441 = " CLK_BASE->S_RDATA_HRDATA[12] = 3.164"
syn_tco442 = " CLK_BASE->S_RDATA_HRDATA[13] = 3.137"
syn_tco443 = " CLK_BASE->S_RDATA_HRDATA[14] = 3.161"
syn_tco444 = " CLK_BASE->S_RDATA_HRDATA[15] = 3.150"
syn_tco445 = " CLK_BASE->S_RDATA_HRDATA[16] = 3.186"
syn_tco446 = " CLK_BASE->S_RDATA_HRDATA[17] = 3.128"
syn_tco447 = " CLK_BASE->S_RDATA_HRDATA[18] = 3.142"
syn_tco448 = " CLK_BASE->S_RDATA_HRDATA[19] = 3.181"
syn_tco449 = " CLK_BASE->S_RDATA_HRDATA[1] = 3.155"
syn_tco450 = " CLK_BASE->S_RDATA_HRDATA[20] = 3.159"
syn_tco451 = " CLK_BASE->S_RDATA_HRDATA[21] = 3.128"
syn_tco452 = " CLK_BASE->S_RDATA_HRDATA[22] = 3.146"
syn_tco453 = " CLK_BASE->S_RDATA_HRDATA[23] = 3.170"
syn_tco454 = " CLK_BASE->S_RDATA_HRDATA[24] = 3.185"
syn_tco455 = " CLK_BASE->S_RDATA_HRDATA[25] = 3.220"
syn_tco456 = " CLK_BASE->S_RDATA_HRDATA[26] = 3.180"
syn_tco457 = " CLK_BASE->S_RDATA_HRDATA[27] = 3.188"
syn_tco458 = " CLK_BASE->S_RDATA_HRDATA[28] = 3.141"
syn_tco459 = " CLK_BASE->S_RDATA_HRDATA[29] = 3.175"
syn_tco460 = " CLK_BASE->S_RDATA_HRDATA[2] = 3.139"
syn_tco461 = " CLK_BASE->S_RDATA_HRDATA[30] = 3.170"
syn_tco462 = " CLK_BASE->S_RDATA_HRDATA[31] = 3.183"
syn_tco463 = " CLK_BASE->S_RDATA_HRDATA[32] = 3.285"
syn_tco464 = " CLK_BASE->S_RDATA_HRDATA[33] = 3.299"
syn_tco465 = " CLK_BASE->S_RDATA_HRDATA[34] = 3.362"
syn_tco466 = " CLK_BASE->S_RDATA_HRDATA[35] = 3.306"
syn_tco467 = " CLK_BASE->S_RDATA_HRDATA[36] = 3.256"
syn_tco468 = " CLK_BASE->S_RDATA_HRDATA[37] = 3.260"
syn_tco469 = " CLK_BASE->S_RDATA_HRDATA[38] = 3.263"
syn_tco470 = " CLK_BASE->S_RDATA_HRDATA[39] = 3.294"
syn_tco471 = " CLK_BASE->S_RDATA_HRDATA[3] = 3.178"
syn_tco472 = " CLK_BASE->S_RDATA_HRDATA[40] = 3.277"
syn_tco473 = " CLK_BASE->S_RDATA_HRDATA[41] = 3.293"
syn_tco474 = " CLK_BASE->S_RDATA_HRDATA[42] = 3.261"
syn_tco475 = " CLK_BASE->S_RDATA_HRDATA[43] = 3.304"
syn_tco476 = " CLK_BASE->S_RDATA_HRDATA[44] = 3.432"
syn_tco477 = " CLK_BASE->S_RDATA_HRDATA[45] = 3.389"
syn_tco478 = " CLK_BASE->S_RDATA_HRDATA[46] = 3.439"
syn_tco479 = " CLK_BASE->S_RDATA_HRDATA[47] = 3.312"
syn_tco480 = " CLK_BASE->S_RDATA_HRDATA[48] = 3.284"
syn_tco481 = " CLK_BASE->S_RDATA_HRDATA[49] = 3.246"
syn_tco482 = " CLK_BASE->S_RDATA_HRDATA[4] = 3.132"
syn_tco483 = " CLK_BASE->S_RDATA_HRDATA[50] = 3.289"
syn_tco484 = " CLK_BASE->S_RDATA_HRDATA[51] = 3.233"
syn_tco485 = " CLK_BASE->S_RDATA_HRDATA[52] = 3.175"
syn_tco486 = " CLK_BASE->S_RDATA_HRDATA[53] = 3.163"
syn_tco487 = " CLK_BASE->S_RDATA_HRDATA[54] = 3.157"
syn_tco488 = " CLK_BASE->S_RDATA_HRDATA[55] = 3.169"
syn_tco489 = " CLK_BASE->S_RDATA_HRDATA[56] = 3.169"
syn_tco490 = " CLK_BASE->S_RDATA_HRDATA[57] = 3.147"
syn_tco491 = " CLK_BASE->S_RDATA_HRDATA[58] = 3.140"
syn_tco492 = " CLK_BASE->S_RDATA_HRDATA[59] = 3.196"
syn_tco493 = " CLK_BASE->S_RDATA_HRDATA[5] = 3.126"
syn_tco494 = " CLK_BASE->S_RDATA_HRDATA[60] = 3.181"
syn_tco495 = " CLK_BASE->S_RDATA_HRDATA[61] = 3.210"
syn_tco496 = " CLK_BASE->S_RDATA_HRDATA[62] = 3.199"
syn_tco497 = " CLK_BASE->S_RDATA_HRDATA[63] = 3.143"
syn_tco498 = " CLK_BASE->S_RDATA_HRDATA[6] = 3.176"
syn_tco499 = " CLK_BASE->S_RDATA_HRDATA[7] = 3.169"
syn_tco500 = " CLK_BASE->S_RDATA_HRDATA[8] = 3.209"
syn_tco501 = " CLK_BASE->S_RDATA_HRDATA[9] = 3.125"
syn_tco502 = " CLK_BASE->S_RID[0] = 3.275"
syn_tco503 = " CLK_BASE->S_RID[1] = 3.215"
syn_tco504 = " CLK_BASE->S_RID[2] = 3.140"
syn_tco505 = " CLK_BASE->S_RID[3] = 3.162"
syn_tco506 = " CLK_BASE->S_RLAST = 3.242"
syn_tco507 = " CLK_BASE->S_RRESP[1] = 3.150"
syn_tco508 = " CLK_BASE->S_RVALID = 3.122"
syn_tco509 = " CLK_BASE->S_WREADY_HREADYOUT = 2.805"
*/
/* synthesis black_box_pad_pin ="RXD3_P,RXD2_P,RXD1_P,RXD0_P,RXD3_N,RXD2_N,RXD1_N,RXD0_N,TXD3_P,TXD2_P,TXD1_P,TXD0_P,TXD3_N,TXD2_N,TXD1_N,TXD0_N" */
output [31:0] APB_PRDATA;
output APB_PREADY;
output APB_PSLVERR;
output [1:0] ATXCLKSTABLE;
output [1:0] EPCS_READY;
output [1:0] EPCS_RXCLK;
output EPCS_RXCLK_0;
output EPCS_RXCLK_1;
output [39:0] EPCS_RXDATA;
output [1:0] EPCS_RXIDLE;
output [1:0] EPCS_RXRSTN;
output [1:0] EPCS_RXVAL;
output [1:0] EPCS_TXCLK;
output EPCS_TXCLK_0;
output EPCS_TXCLK_1;
output [1:0] EPCS_TXRSTN;
output FATC_RESET_N;
output H2FCALIB0;
output H2FCALIB1;
output [31:0] M2_ARADDR;
output [1:0] M2_ARBURST;
output [3:0] M2_ARID;
output [3:0] M2_ARLEN;
output [1:0] M2_ARSIZE;
output M2_ARVALID;
output [31:0] M2_AWADDR_HADDR;
output [1:0] M2_AWBURST_HTRANS;
output [3:0] M2_AWID;
output [3:0] M2_AWLEN_HBURST;
output [1:0] M2_AWSIZE_HSIZE;
output M2_AWVALID_HWRITE;
output M2_BREADY;
output M2_RREADY;
output [63:0] M2_WDATA_HWDATA;
output [3:0] M2_WID;
output M2_WLAST;
output [7:0] M2_WSTRB;
output M2_WVALID;
output [31:0] M_ARADDR;
output [1:0] M_ARBURST;
output [3:0] M_ARID;
output [3:0] M_ARLEN;
output [1:0] M_ARSIZE;
output M_ARVALID;
output [31:0] M_AWADDR_HADDR;
output [1:0] M_AWBURST_HTRANS;
output [3:0] M_AWID;
output [3:0] M_AWLEN_HBURST;
output [1:0] M_AWSIZE_HSIZE;
output M_AWVALID_HWRITE;
output M_BREADY;
output M_RREADY;
output [63:0] M_WDATA_HWDATA;
output [3:0] M_WID;
output M_WLAST;
output [7:0] M_WSTRB;
output M_WVALID;
output [5:0] PCIE2_LTSSM;
output PCIE2_SYSTEM_INT;
output PCIE2_WAKE_N;
output [5:0] PCIE_LTSSM;
output PCIE_SYSTEM_INT;
output PLL_LOCK_INT;
output PLL_LOCKLOST_INT;
output S2_ARREADY;
output S2_AWREADY;
output [3:0] S2_BID;
output [1:0] S2_BRESP_HRESP;
output S2_BVALID;
output [63:0] S2_RDATA_HRDATA;
output [3:0] S2_RID;
output S2_RLAST;
output [1:0] S2_RRESP;
output S2_RVALID;
output S2_WREADY_HREADYOUT;
output S_ARREADY;
output S_AWREADY;
output [3:0] S_BID;
output [1:0] S_BRESP_HRESP;
output S_BVALID;
output [63:0] S_RDATA_HRDATA;
output [3:0] S_RID;
output S_RLAST;
output [1:0] S_RRESP;
output S_RVALID;
output S_WREADY_HREADYOUT;
output SPLL_LOCK;
output WAKE_N;
output XAUI_OUT_CLK;
input  APB_CLK;
input  [14:2] APB_PADDR;
input  APB_PENABLE;
input  APB_PSEL;
input  [31:0] APB_PWDATA;
input  APB_PWRITE;
input  APB_RSTN;
input  CLK_BASE;
input  [1:0] EPCS_PWRDN;
input  [1:0] EPCS_RSTN;
input  [1:0] EPCS_RXERR;
input  [39:0] EPCS_TXDATA;
input  [1:0] EPCS_TXOOB;
input  [1:0] EPCS_TXVAL;
input  F2HCALIB0;
input  F2HCALIB1;
input  FAB_PLL_LOCK;
input  FAB_REF_CLK;
input  M2_ARREADY;
input  M2_AWREADY;
input  [3:0] M2_BID;
input  [1:0] M2_BRESP_HRESP;
input  M2_BVALID;
input  [63:0] M2_RDATA_HRDATA;
input  [3:0] M2_RID;
input  M2_RLAST;
input  [1:0] M2_RRESP;
input  M2_RVALID;
input  M2_WREADY_HREADY;
input  M_ARREADY;
input  M_AWREADY;
input  [3:0] M_BID;
input  [1:0] M_BRESP_HRESP;
input  M_BVALID;
input  [63:0] M_RDATA_HRDATA;
input  [3:0] M_RID;
input  M_RLAST;
input  [1:0] M_RRESP;
input  M_RVALID;
input  M_WREADY_HREADY;
input  [3:0] PCIE2_INTERRUPT;
input  PCIE2_PERST_N;
input  PCIE2_SERDESIF_CORE_RESET_N;
input  PCIE2_WAKE_REQ;
input  [3:0] PCIE_INTERRUPT;
input  PERST_N;
input  [31:0] S2_ARADDR;
input  [1:0] S2_ARBURST;
input  [3:0] S2_ARID;
input  [3:0] S2_ARLEN;
input  [1:0] S2_ARLOCK;
input  [1:0] S2_ARSIZE;
input  S2_ARVALID;
input  [31:0] S2_AWADDR_HADDR;
input  [1:0] S2_AWBURST_HTRANS;
input  [3:0] S2_AWID_HSEL;
input  [3:0] S2_AWLEN_HBURST;
input  [1:0] S2_AWLOCK;
input  [1:0] S2_AWSIZE_HSIZE;
input  S2_AWVALID_HWRITE;
input  S2_BREADY_HREADY;
input  S2_RREADY;
input  [63:0] S2_WDATA_HWDATA;
input  [3:0] S2_WID;
input  S2_WLAST;
input  [7:0] S2_WSTRB;
input  S2_WVALID;
input  [31:0] S_ARADDR;
input  [1:0] S_ARBURST;
input  [3:0] S_ARID;
input  [3:0] S_ARLEN;
input  [1:0] S_ARLOCK;
input  [1:0] S_ARSIZE;
input  S_ARVALID;
input  [31:0] S_AWADDR_HADDR;
input  [1:0] S_AWBURST_HTRANS;
input  [3:0] S_AWID_HSEL;
input  [3:0] S_AWLEN_HBURST;
input  [1:0] S_AWLOCK;
input  [1:0] S_AWSIZE_HSIZE;
input  S_AWVALID_HWRITE;
input  S_BREADY_HREADY;
input  S_RREADY;
input  [63:0] S_WDATA_HWDATA;
input  [3:0] S_WID;
input  S_WLAST;
input  [7:0] S_WSTRB;
input  S_WVALID;
input  SERDESIF_CORE_RESET_N;
input  SERDESIF_PHY_RESET_N;
input  WAKE_REQ;
input  XAUI_FB_CLK;
input  RXD3_P;
input  RXD2_P;
input  RXD1_P;
input  RXD0_P;
input  RXD3_N;
input  RXD2_N;
input  RXD1_N;
input  RXD0_N;
output TXD3_P;
output TXD2_P;
output TXD1_P;
output TXD0_P;
output TXD3_N;
output TXD2_N;
output TXD1_N;
output TXD0_N;
input  REFCLK0;
input  REFCLK1;
parameter INIT = 'h0;
parameter ACT_CONFIG = "";
parameter ACT_SIM = 0;

endmodule
