`timescale 1 ns/100 ps
// Version: 


module SERDESIF_075(
       APB_PRDATA,
       APB_PREADY,
       APB_PSLVERR,
       ATXCLKSTABLE,
       EPCS_READY,
       EPCS_RXCLK,
       EPCS_RXCLK_0,
       EPCS_RXCLK_1,
       EPCS_RXDATA,
       EPCS_RXIDLE,
       EPCS_RXRSTN,
       EPCS_RXVAL,
       EPCS_TXCLK,
       EPCS_TXCLK_0,
       EPCS_TXCLK_1,
       EPCS_TXRSTN,
       FATC_RESET_N,
       H2FCALIB0,
       H2FCALIB1,
       M2_ARADDR,
       M2_ARBURST,
       M2_ARID,
       M2_ARLEN,
       M2_ARSIZE,
       M2_ARVALID,
       M2_AWADDR_HADDR,
       M2_AWBURST_HTRANS,
       M2_AWID,
       M2_AWLEN_HBURST,
       M2_AWSIZE_HSIZE,
       M2_AWVALID_HWRITE,
       M2_BREADY,
       M2_RREADY,
       M2_WDATA_HWDATA,
       M2_WID,
       M2_WLAST,
       M2_WSTRB,
       M2_WVALID,
       M_ARADDR,
       M_ARBURST,
       M_ARID,
       M_ARLEN,
       M_ARSIZE,
       M_ARVALID,
       M_AWADDR_HADDR,
       M_AWBURST_HTRANS,
       M_AWID,
       M_AWLEN_HBURST,
       M_AWSIZE_HSIZE,
       M_AWVALID_HWRITE,
       M_BREADY,
       M_RREADY,
       M_WDATA_HWDATA,
       M_WID,
       M_WLAST,
       M_WSTRB,
       M_WVALID,
       PCIE2_LTSSM,
       PCIE2_SYSTEM_INT,
       PCIE2_WAKE_N,
       PCIE_LTSSM,
       PCIE_SYSTEM_INT,
       PLL_LOCK_INT,
       PLL_LOCKLOST_INT,
       S2_ARREADY,
       S2_AWREADY,
       S2_BID,
       S2_BRESP_HRESP,
       S2_BVALID,
       S2_RDATA_HRDATA,
       S2_RID,
       S2_RLAST,
       S2_RRESP,
       S2_RVALID,
       S2_WREADY_HREADYOUT,
       S_ARREADY,
       S_AWREADY,
       S_BID,
       S_BRESP_HRESP,
       S_BVALID,
       S_RDATA_HRDATA,
       S_RID,
       S_RLAST,
       S_RRESP,
       S_RVALID,
       S_WREADY_HREADYOUT,
       SPLL_LOCK,
       WAKE_N,
       XAUI_OUT_CLK,
       APB_CLK,
       APB_PADDR,
       APB_PENABLE,
       APB_PSEL,
       APB_PWDATA,
       APB_PWRITE,
       APB_RSTN,
       CLK_BASE,
       EPCS_PWRDN,
       EPCS_RSTN,
       EPCS_RXERR,
       EPCS_TXDATA,
       EPCS_TXOOB,
       EPCS_TXVAL,
       F2HCALIB0,
       F2HCALIB1,
       FAB_PLL_LOCK,
       FAB_REF_CLK,
       M2_ARREADY,
       M2_AWREADY,
       M2_BID,
       M2_BRESP_HRESP,
       M2_BVALID,
       M2_RDATA_HRDATA,
       M2_RID,
       M2_RLAST,
       M2_RRESP,
       M2_RVALID,
       M2_WREADY_HREADY,
       M_ARREADY,
       M_AWREADY,
       M_BID,
       M_BRESP_HRESP,
       M_BVALID,
       M_RDATA_HRDATA,
       M_RID,
       M_RLAST,
       M_RRESP,
       M_RVALID,
       M_WREADY_HREADY,
       PCIE2_INTERRUPT,
       PCIE2_PERST_N,
       PCIE2_SERDESIF_CORE_RESET_N,
       PCIE2_WAKE_REQ,
       PCIE_INTERRUPT,
       PERST_N,
       S2_ARADDR,
       S2_ARBURST,
       S2_ARID,
       S2_ARLEN,
       S2_ARLOCK,
       S2_ARSIZE,
       S2_ARVALID,
       S2_AWADDR_HADDR,
       S2_AWBURST_HTRANS,
       S2_AWID_HSEL,
       S2_AWLEN_HBURST,
       S2_AWLOCK,
       S2_AWSIZE_HSIZE,
       S2_AWVALID_HWRITE,
       S2_BREADY_HREADY,
       S2_RREADY,
       S2_WDATA_HWDATA,
       S2_WID,
       S2_WLAST,
       S2_WSTRB,
       S2_WVALID,
       S_ARADDR,
       S_ARBURST,
       S_ARID,
       S_ARLEN,
       S_ARLOCK,
       S_ARSIZE,
       S_ARVALID,
       S_AWADDR_HADDR,
       S_AWBURST_HTRANS,
       S_AWID_HSEL,
       S_AWLEN_HBURST,
       S_AWLOCK,
       S_AWSIZE_HSIZE,
       S_AWVALID_HWRITE,
       S_BREADY_HREADY,
       S_RREADY,
       S_WDATA_HWDATA,
       S_WID,
       S_WLAST,
       S_WSTRB,
       S_WVALID,
       SERDESIF_CORE_RESET_N,
       SERDESIF_PHY_RESET_N,
       WAKE_REQ,
       XAUI_FB_CLK,
       RXD3_P,
       RXD2_P,
       RXD1_P,
       RXD0_P,
       RXD3_N,
       RXD2_N,
       RXD1_N,
       RXD0_N,
       TXD3_P,
       TXD2_P,
       TXD1_P,
       TXD0_P,
       TXD3_N,
       TXD2_N,
       TXD1_N,
       TXD0_N,
       REFCLK0,
       REFCLK1
    )
/* synthesis black_box

pragma attribute SERDESIF_075 ment_tsu0 APB_PADDR[10]->APB_CLK+3.791
pragma attribute SERDESIF_075 ment_tsu1 APB_PADDR[11]->APB_CLK+3.498
pragma attribute SERDESIF_075 ment_tsu2 APB_PADDR[12]->APB_CLK+3.309
pragma attribute SERDESIF_075 ment_tsu3 APB_PADDR[13]->APB_CLK+3.076
pragma attribute SERDESIF_075 ment_tsu4 APB_PADDR[14]->APB_CLK+2.521
pragma attribute SERDESIF_075 ment_tsu5 APB_PADDR[2]->APB_CLK+2.929
pragma attribute SERDESIF_075 ment_tsu6 APB_PADDR[3]->APB_CLK+3.244
pragma attribute SERDESIF_075 ment_tsu7 APB_PADDR[4]->APB_CLK+2.893
pragma attribute SERDESIF_075 ment_tsu8 APB_PADDR[5]->APB_CLK+3.290
pragma attribute SERDESIF_075 ment_tsu9 APB_PADDR[6]->APB_CLK+2.853
pragma attribute SERDESIF_075 ment_tsu10 APB_PADDR[7]->APB_CLK+2.851
pragma attribute SERDESIF_075 ment_tsu11 APB_PADDR[8]->APB_CLK+3.480
pragma attribute SERDESIF_075 ment_tsu12 APB_PADDR[9]->APB_CLK+3.473
pragma attribute SERDESIF_075 ment_tsu13 APB_PENABLE->APB_CLK+0.833
pragma attribute SERDESIF_075 ment_tsu14 APB_PSEL->APB_CLK+2.830
pragma attribute SERDESIF_075 ment_tsu15 APB_PWDATA[0]->APB_CLK+1.294
pragma attribute SERDESIF_075 ment_tsu16 APB_PWDATA[10]->APB_CLK+0.494
pragma attribute SERDESIF_075 ment_tsu17 APB_PWDATA[11]->APB_CLK+0.581
pragma attribute SERDESIF_075 ment_tsu18 APB_PWDATA[12]->APB_CLK+0.831
pragma attribute SERDESIF_075 ment_tsu19 APB_PWDATA[13]->APB_CLK+0.725
pragma attribute SERDESIF_075 ment_tsu20 APB_PWDATA[14]->APB_CLK+0.897
pragma attribute SERDESIF_075 ment_tsu21 APB_PWDATA[15]->APB_CLK+0.713
pragma attribute SERDESIF_075 ment_tsu22 APB_PWDATA[16]->APB_CLK+0.813
pragma attribute SERDESIF_075 ment_tsu23 APB_PWDATA[17]->APB_CLK+0.747
pragma attribute SERDESIF_075 ment_tsu24 APB_PWDATA[18]->APB_CLK+0.748
pragma attribute SERDESIF_075 ment_tsu25 APB_PWDATA[19]->APB_CLK+0.954
pragma attribute SERDESIF_075 ment_tsu26 APB_PWDATA[1]->APB_CLK+1.879
pragma attribute SERDESIF_075 ment_tsu27 APB_PWDATA[20]->APB_CLK+0.803
pragma attribute SERDESIF_075 ment_tsu28 APB_PWDATA[21]->APB_CLK+0.460
pragma attribute SERDESIF_075 ment_tsu29 APB_PWDATA[22]->APB_CLK+0.516
pragma attribute SERDESIF_075 ment_tsu30 APB_PWDATA[23]->APB_CLK+0.496
pragma attribute SERDESIF_075 ment_tsu31 APB_PWDATA[24]->APB_CLK+0.642
pragma attribute SERDESIF_075 ment_tsu32 APB_PWDATA[25]->APB_CLK+0.509
pragma attribute SERDESIF_075 ment_tsu33 APB_PWDATA[26]->APB_CLK+0.421
pragma attribute SERDESIF_075 ment_tsu34 APB_PWDATA[27]->APB_CLK+0.546
pragma attribute SERDESIF_075 ment_tsu35 APB_PWDATA[28]->APB_CLK+0.087
pragma attribute SERDESIF_075 ment_tsu36 APB_PWDATA[29]->APB_CLK+-0.005
pragma attribute SERDESIF_075 ment_tsu37 APB_PWDATA[2]->APB_CLK+1.743
pragma attribute SERDESIF_075 ment_tsu38 APB_PWDATA[30]->APB_CLK+0.556
pragma attribute SERDESIF_075 ment_tsu39 APB_PWDATA[31]->APB_CLK+0.054
pragma attribute SERDESIF_075 ment_tsu40 APB_PWDATA[3]->APB_CLK+1.950
pragma attribute SERDESIF_075 ment_tsu41 APB_PWDATA[4]->APB_CLK+1.925
pragma attribute SERDESIF_075 ment_tsu42 APB_PWDATA[5]->APB_CLK+1.226
pragma attribute SERDESIF_075 ment_tsu43 APB_PWDATA[6]->APB_CLK+1.954
pragma attribute SERDESIF_075 ment_tsu44 APB_PWDATA[7]->APB_CLK+0.928
pragma attribute SERDESIF_075 ment_tsu45 APB_PWDATA[8]->APB_CLK+0.693
pragma attribute SERDESIF_075 ment_tsu46 APB_PWDATA[9]->APB_CLK+0.849
pragma attribute SERDESIF_075 ment_tsu47 APB_PWRITE->APB_CLK+1.751
pragma attribute SERDESIF_075 ment_tsu48 M2_ARREADY->CLK_BASE+0.920
pragma attribute SERDESIF_075 ment_tsu49 M2_AWREADY->CLK_BASE+0.812
pragma attribute SERDESIF_075 ment_tsu50 M2_BID[0]->CLK_BASE+0.079
pragma attribute SERDESIF_075 ment_tsu51 M2_BRESP_HRESP[0]->CLK_BASE+0.119
pragma attribute SERDESIF_075 ment_tsu52 M2_BVALID->CLK_BASE+0.892
pragma attribute SERDESIF_075 ment_tsu53 M2_RDATA_HRDATA[0]->CLK_BASE+0.632
pragma attribute SERDESIF_075 ment_tsu54 M2_RDATA_HRDATA[10]->CLK_BASE+0.666
pragma attribute SERDESIF_075 ment_tsu55 M2_RDATA_HRDATA[11]->CLK_BASE+0.530
pragma attribute SERDESIF_075 ment_tsu56 M2_RDATA_HRDATA[12]->CLK_BASE+0.706
pragma attribute SERDESIF_075 ment_tsu57 M2_RDATA_HRDATA[13]->CLK_BASE+0.283
pragma attribute SERDESIF_075 ment_tsu58 M2_RDATA_HRDATA[14]->CLK_BASE+0.626
pragma attribute SERDESIF_075 ment_tsu59 M2_RDATA_HRDATA[15]->CLK_BASE+0.499
pragma attribute SERDESIF_075 ment_tsu60 M2_RDATA_HRDATA[16]->CLK_BASE+0.761
pragma attribute SERDESIF_075 ment_tsu61 M2_RDATA_HRDATA[17]->CLK_BASE+0.529
pragma attribute SERDESIF_075 ment_tsu62 M2_RDATA_HRDATA[18]->CLK_BASE+0.721
pragma attribute SERDESIF_075 ment_tsu63 M2_RDATA_HRDATA[19]->CLK_BASE+0.751
pragma attribute SERDESIF_075 ment_tsu64 M2_RDATA_HRDATA[1]->CLK_BASE+0.691
pragma attribute SERDESIF_075 ment_tsu65 M2_RDATA_HRDATA[20]->CLK_BASE+0.417
pragma attribute SERDESIF_075 ment_tsu66 M2_RDATA_HRDATA[21]->CLK_BASE+0.449
pragma attribute SERDESIF_075 ment_tsu67 M2_RDATA_HRDATA[22]->CLK_BASE+0.280
pragma attribute SERDESIF_075 ment_tsu68 M2_RDATA_HRDATA[23]->CLK_BASE+0.657
pragma attribute SERDESIF_075 ment_tsu69 M2_RDATA_HRDATA[24]->CLK_BASE+0.750
pragma attribute SERDESIF_075 ment_tsu70 M2_RDATA_HRDATA[25]->CLK_BASE+0.841
pragma attribute SERDESIF_075 ment_tsu71 M2_RDATA_HRDATA[26]->CLK_BASE+0.572
pragma attribute SERDESIF_075 ment_tsu72 M2_RDATA_HRDATA[27]->CLK_BASE+0.174
pragma attribute SERDESIF_075 ment_tsu73 M2_RDATA_HRDATA[28]->CLK_BASE+0.712
pragma attribute SERDESIF_075 ment_tsu74 M2_RDATA_HRDATA[29]->CLK_BASE+0.707
pragma attribute SERDESIF_075 ment_tsu75 M2_RDATA_HRDATA[2]->CLK_BASE+0.769
pragma attribute SERDESIF_075 ment_tsu76 M2_RDATA_HRDATA[30]->CLK_BASE+0.389
pragma attribute SERDESIF_075 ment_tsu77 M2_RDATA_HRDATA[31]->CLK_BASE+0.729
pragma attribute SERDESIF_075 ment_tsu78 M2_RDATA_HRDATA[32]->CLK_BASE+0.879
pragma attribute SERDESIF_075 ment_tsu79 M2_RDATA_HRDATA[33]->CLK_BASE+0.853
pragma attribute SERDESIF_075 ment_tsu80 M2_RDATA_HRDATA[34]->CLK_BASE+-0.003
pragma attribute SERDESIF_075 ment_tsu81 M2_RDATA_HRDATA[35]->CLK_BASE+0.191
pragma attribute SERDESIF_075 ment_tsu82 M2_RDATA_HRDATA[36]->CLK_BASE+0.532
pragma attribute SERDESIF_075 ment_tsu83 M2_RDATA_HRDATA[37]->CLK_BASE+0.525
pragma attribute SERDESIF_075 ment_tsu84 M2_RDATA_HRDATA[38]->CLK_BASE+0.953
pragma attribute SERDESIF_075 ment_tsu85 M2_RDATA_HRDATA[39]->CLK_BASE+0.458
pragma attribute SERDESIF_075 ment_tsu86 M2_RDATA_HRDATA[3]->CLK_BASE+0.830
pragma attribute SERDESIF_075 ment_tsu87 M2_RDATA_HRDATA[40]->CLK_BASE+0.557
pragma attribute SERDESIF_075 ment_tsu88 M2_RDATA_HRDATA[41]->CLK_BASE+0.571
pragma attribute SERDESIF_075 ment_tsu89 M2_RDATA_HRDATA[42]->CLK_BASE+0.379
pragma attribute SERDESIF_075 ment_tsu90 M2_RDATA_HRDATA[43]->CLK_BASE+0.795
pragma attribute SERDESIF_075 ment_tsu91 M2_RDATA_HRDATA[44]->CLK_BASE+0.942
pragma attribute SERDESIF_075 ment_tsu92 M2_RDATA_HRDATA[45]->CLK_BASE+0.537
pragma attribute SERDESIF_075 ment_tsu93 M2_RDATA_HRDATA[46]->CLK_BASE+0.791
pragma attribute SERDESIF_075 ment_tsu94 M2_RDATA_HRDATA[47]->CLK_BASE+0.021
pragma attribute SERDESIF_075 ment_tsu95 M2_RDATA_HRDATA[48]->CLK_BASE+0.436
pragma attribute SERDESIF_075 ment_tsu96 M2_RDATA_HRDATA[49]->CLK_BASE+0.803
pragma attribute SERDESIF_075 ment_tsu97 M2_RDATA_HRDATA[4]->CLK_BASE+0.530
pragma attribute SERDESIF_075 ment_tsu98 M2_RDATA_HRDATA[50]->CLK_BASE+0.186
pragma attribute SERDESIF_075 ment_tsu99 M2_RDATA_HRDATA[51]->CLK_BASE+0.894
pragma attribute SERDESIF_075 ment_tsu100 M2_RDATA_HRDATA[52]->CLK_BASE+0.495
pragma attribute SERDESIF_075 ment_tsu101 M2_RDATA_HRDATA[53]->CLK_BASE+0.649
pragma attribute SERDESIF_075 ment_tsu102 M2_RDATA_HRDATA[54]->CLK_BASE+0.518
pragma attribute SERDESIF_075 ment_tsu103 M2_RDATA_HRDATA[55]->CLK_BASE+0.620
pragma attribute SERDESIF_075 ment_tsu104 M2_RDATA_HRDATA[56]->CLK_BASE+0.717
pragma attribute SERDESIF_075 ment_tsu105 M2_RDATA_HRDATA[57]->CLK_BASE+0.690
pragma attribute SERDESIF_075 ment_tsu106 M2_RDATA_HRDATA[58]->CLK_BASE+0.589
pragma attribute SERDESIF_075 ment_tsu107 M2_RDATA_HRDATA[59]->CLK_BASE+0.927
pragma attribute SERDESIF_075 ment_tsu108 M2_RDATA_HRDATA[5]->CLK_BASE+0.580
pragma attribute SERDESIF_075 ment_tsu109 M2_RDATA_HRDATA[60]->CLK_BASE+0.524
pragma attribute SERDESIF_075 ment_tsu110 M2_RDATA_HRDATA[61]->CLK_BASE+0.329
pragma attribute SERDESIF_075 ment_tsu111 M2_RDATA_HRDATA[62]->CLK_BASE+0.598
pragma attribute SERDESIF_075 ment_tsu112 M2_RDATA_HRDATA[63]->CLK_BASE+0.822
pragma attribute SERDESIF_075 ment_tsu113 M2_RDATA_HRDATA[6]->CLK_BASE+0.806
pragma attribute SERDESIF_075 ment_tsu114 M2_RDATA_HRDATA[7]->CLK_BASE+0.747
pragma attribute SERDESIF_075 ment_tsu115 M2_RDATA_HRDATA[8]->CLK_BASE+0.325
pragma attribute SERDESIF_075 ment_tsu116 M2_RDATA_HRDATA[9]->CLK_BASE+0.655
pragma attribute SERDESIF_075 ment_tsu117 M2_RID[0]->CLK_BASE+0.600
pragma attribute SERDESIF_075 ment_tsu118 M2_RID[1]->CLK_BASE+0.634
pragma attribute SERDESIF_075 ment_tsu119 M2_RID[2]->CLK_BASE+0.103
pragma attribute SERDESIF_075 ment_tsu120 M2_RID[3]->CLK_BASE+0.533
pragma attribute SERDESIF_075 ment_tsu121 M2_RLAST->CLK_BASE+0.628
pragma attribute SERDESIF_075 ment_tsu122 M2_RRESP[0]->CLK_BASE+0.216
pragma attribute SERDESIF_075 ment_tsu123 M2_RRESP[1]->CLK_BASE+0.721
pragma attribute SERDESIF_075 ment_tsu124 M2_RVALID->CLK_BASE+0.936
pragma attribute SERDESIF_075 ment_tsu125 M2_WREADY_HREADY->CLK_BASE+0.991
pragma attribute SERDESIF_075 ment_tsu126 M_ARREADY->CLK_BASE+0.860
pragma attribute SERDESIF_075 ment_tsu127 M_AWREADY->CLK_BASE+1.008
pragma attribute SERDESIF_075 ment_tsu128 M_BID[0]->CLK_BASE+0.564
pragma attribute SERDESIF_075 ment_tsu129 M_BRESP_HRESP[0]->CLK_BASE+0.392
pragma attribute SERDESIF_075 ment_tsu130 M_BVALID->CLK_BASE+0.596
pragma attribute SERDESIF_075 ment_tsu131 M_RDATA_HRDATA[0]->CLK_BASE+0.787
pragma attribute SERDESIF_075 ment_tsu132 M_RDATA_HRDATA[10]->CLK_BASE+0.781
pragma attribute SERDESIF_075 ment_tsu133 M_RDATA_HRDATA[11]->CLK_BASE+0.977
pragma attribute SERDESIF_075 ment_tsu134 M_RDATA_HRDATA[12]->CLK_BASE+0.553
pragma attribute SERDESIF_075 ment_tsu135 M_RDATA_HRDATA[13]->CLK_BASE+0.804
pragma attribute SERDESIF_075 ment_tsu136 M_RDATA_HRDATA[14]->CLK_BASE+0.605
pragma attribute SERDESIF_075 ment_tsu137 M_RDATA_HRDATA[15]->CLK_BASE+0.914
pragma attribute SERDESIF_075 ment_tsu138 M_RDATA_HRDATA[16]->CLK_BASE+0.670
pragma attribute SERDESIF_075 ment_tsu139 M_RDATA_HRDATA[17]->CLK_BASE+0.579
pragma attribute SERDESIF_075 ment_tsu140 M_RDATA_HRDATA[18]->CLK_BASE+0.557
pragma attribute SERDESIF_075 ment_tsu141 M_RDATA_HRDATA[19]->CLK_BASE+0.732
pragma attribute SERDESIF_075 ment_tsu142 M_RDATA_HRDATA[1]->CLK_BASE+0.748
pragma attribute SERDESIF_075 ment_tsu143 M_RDATA_HRDATA[20]->CLK_BASE+0.604
pragma attribute SERDESIF_075 ment_tsu144 M_RDATA_HRDATA[21]->CLK_BASE+0.795
pragma attribute SERDESIF_075 ment_tsu145 M_RDATA_HRDATA[22]->CLK_BASE+0.960
pragma attribute SERDESIF_075 ment_tsu146 M_RDATA_HRDATA[23]->CLK_BASE+0.900
pragma attribute SERDESIF_075 ment_tsu147 M_RDATA_HRDATA[24]->CLK_BASE+0.339
pragma attribute SERDESIF_075 ment_tsu148 M_RDATA_HRDATA[25]->CLK_BASE+0.755
pragma attribute SERDESIF_075 ment_tsu149 M_RDATA_HRDATA[26]->CLK_BASE+0.537
pragma attribute SERDESIF_075 ment_tsu150 M_RDATA_HRDATA[27]->CLK_BASE+0.600
pragma attribute SERDESIF_075 ment_tsu151 M_RDATA_HRDATA[28]->CLK_BASE+0.771
pragma attribute SERDESIF_075 ment_tsu152 M_RDATA_HRDATA[29]->CLK_BASE+0.531
pragma attribute SERDESIF_075 ment_tsu153 M_RDATA_HRDATA[2]->CLK_BASE+0.934
pragma attribute SERDESIF_075 ment_tsu154 M_RDATA_HRDATA[30]->CLK_BASE+0.567
pragma attribute SERDESIF_075 ment_tsu155 M_RDATA_HRDATA[31]->CLK_BASE+0.631
pragma attribute SERDESIF_075 ment_tsu156 M_RDATA_HRDATA[32]->CLK_BASE+0.737
pragma attribute SERDESIF_075 ment_tsu157 M_RDATA_HRDATA[33]->CLK_BASE+0.538
pragma attribute SERDESIF_075 ment_tsu158 M_RDATA_HRDATA[34]->CLK_BASE+0.756
pragma attribute SERDESIF_075 ment_tsu159 M_RDATA_HRDATA[35]->CLK_BASE+0.628
pragma attribute SERDESIF_075 ment_tsu160 M_RDATA_HRDATA[36]->CLK_BASE+0.282
pragma attribute SERDESIF_075 ment_tsu161 M_RDATA_HRDATA[37]->CLK_BASE+0.847
pragma attribute SERDESIF_075 ment_tsu162 M_RDATA_HRDATA[38]->CLK_BASE+0.689
pragma attribute SERDESIF_075 ment_tsu163 M_RDATA_HRDATA[39]->CLK_BASE+0.941
pragma attribute SERDESIF_075 ment_tsu164 M_RDATA_HRDATA[3]->CLK_BASE+0.868
pragma attribute SERDESIF_075 ment_tsu165 M_RDATA_HRDATA[40]->CLK_BASE+0.700
pragma attribute SERDESIF_075 ment_tsu166 M_RDATA_HRDATA[41]->CLK_BASE+0.798
pragma attribute SERDESIF_075 ment_tsu167 M_RDATA_HRDATA[42]->CLK_BASE+0.902
pragma attribute SERDESIF_075 ment_tsu168 M_RDATA_HRDATA[43]->CLK_BASE+0.707
pragma attribute SERDESIF_075 ment_tsu169 M_RDATA_HRDATA[44]->CLK_BASE+0.877
pragma attribute SERDESIF_075 ment_tsu170 M_RDATA_HRDATA[45]->CLK_BASE+0.595
pragma attribute SERDESIF_075 ment_tsu171 M_RDATA_HRDATA[46]->CLK_BASE+0.929
pragma attribute SERDESIF_075 ment_tsu172 M_RDATA_HRDATA[47]->CLK_BASE+0.827
pragma attribute SERDESIF_075 ment_tsu173 M_RDATA_HRDATA[48]->CLK_BASE+0.532
pragma attribute SERDESIF_075 ment_tsu174 M_RDATA_HRDATA[49]->CLK_BASE+0.801
pragma attribute SERDESIF_075 ment_tsu175 M_RDATA_HRDATA[4]->CLK_BASE+0.734
pragma attribute SERDESIF_075 ment_tsu176 M_RDATA_HRDATA[50]->CLK_BASE+0.835
pragma attribute SERDESIF_075 ment_tsu177 M_RDATA_HRDATA[51]->CLK_BASE+0.887
pragma attribute SERDESIF_075 ment_tsu178 M_RDATA_HRDATA[52]->CLK_BASE+0.889
pragma attribute SERDESIF_075 ment_tsu179 M_RDATA_HRDATA[53]->CLK_BASE+0.745
pragma attribute SERDESIF_075 ment_tsu180 M_RDATA_HRDATA[54]->CLK_BASE+0.768
pragma attribute SERDESIF_075 ment_tsu181 M_RDATA_HRDATA[55]->CLK_BASE+0.607
pragma attribute SERDESIF_075 ment_tsu182 M_RDATA_HRDATA[56]->CLK_BASE+0.820
pragma attribute SERDESIF_075 ment_tsu183 M_RDATA_HRDATA[57]->CLK_BASE+0.295
pragma attribute SERDESIF_075 ment_tsu184 M_RDATA_HRDATA[58]->CLK_BASE+0.414
pragma attribute SERDESIF_075 ment_tsu185 M_RDATA_HRDATA[59]->CLK_BASE+0.920
pragma attribute SERDESIF_075 ment_tsu186 M_RDATA_HRDATA[5]->CLK_BASE+0.852
pragma attribute SERDESIF_075 ment_tsu187 M_RDATA_HRDATA[60]->CLK_BASE+0.448
pragma attribute SERDESIF_075 ment_tsu188 M_RDATA_HRDATA[61]->CLK_BASE+0.785
pragma attribute SERDESIF_075 ment_tsu189 M_RDATA_HRDATA[62]->CLK_BASE+0.458
pragma attribute SERDESIF_075 ment_tsu190 M_RDATA_HRDATA[63]->CLK_BASE+0.884
pragma attribute SERDESIF_075 ment_tsu191 M_RDATA_HRDATA[6]->CLK_BASE+0.401
pragma attribute SERDESIF_075 ment_tsu192 M_RDATA_HRDATA[7]->CLK_BASE+0.623
pragma attribute SERDESIF_075 ment_tsu193 M_RDATA_HRDATA[8]->CLK_BASE+0.911
pragma attribute SERDESIF_075 ment_tsu194 M_RDATA_HRDATA[9]->CLK_BASE+0.709
pragma attribute SERDESIF_075 ment_tsu195 M_RID[0]->CLK_BASE+0.596
pragma attribute SERDESIF_075 ment_tsu196 M_RID[1]->CLK_BASE+0.114
pragma attribute SERDESIF_075 ment_tsu197 M_RID[2]->CLK_BASE+0.661
pragma attribute SERDESIF_075 ment_tsu198 M_RID[3]->CLK_BASE+0.561
pragma attribute SERDESIF_075 ment_tsu199 M_RLAST->CLK_BASE+0.791
pragma attribute SERDESIF_075 ment_tsu200 M_RRESP[0]->CLK_BASE+0.741
pragma attribute SERDESIF_075 ment_tsu201 M_RRESP[1]->CLK_BASE+0.530
pragma attribute SERDESIF_075 ment_tsu202 M_RVALID->CLK_BASE+0.348
pragma attribute SERDESIF_075 ment_tsu203 M_WREADY_HREADY->CLK_BASE+1.052
pragma attribute SERDESIF_075 ment_tsu204 S2_ARADDR[0]->CLK_BASE+0.564
pragma attribute SERDESIF_075 ment_tsu205 S2_ARADDR[10]->CLK_BASE+0.454
pragma attribute SERDESIF_075 ment_tsu206 S2_ARADDR[11]->CLK_BASE+0.669
pragma attribute SERDESIF_075 ment_tsu207 S2_ARADDR[12]->CLK_BASE+0.169
pragma attribute SERDESIF_075 ment_tsu208 S2_ARADDR[13]->CLK_BASE+0.143
pragma attribute SERDESIF_075 ment_tsu209 S2_ARADDR[14]->CLK_BASE+0.487
pragma attribute SERDESIF_075 ment_tsu210 S2_ARADDR[15]->CLK_BASE+0.468
pragma attribute SERDESIF_075 ment_tsu211 S2_ARADDR[16]->CLK_BASE+0.135
pragma attribute SERDESIF_075 ment_tsu212 S2_ARADDR[17]->CLK_BASE+0.110
pragma attribute SERDESIF_075 ment_tsu213 S2_ARADDR[18]->CLK_BASE+0.972
pragma attribute SERDESIF_075 ment_tsu214 S2_ARADDR[19]->CLK_BASE+0.432
pragma attribute SERDESIF_075 ment_tsu215 S2_ARADDR[1]->CLK_BASE+0.552
pragma attribute SERDESIF_075 ment_tsu216 S2_ARADDR[20]->CLK_BASE+0.414
pragma attribute SERDESIF_075 ment_tsu217 S2_ARADDR[21]->CLK_BASE+0.431
pragma attribute SERDESIF_075 ment_tsu218 S2_ARADDR[22]->CLK_BASE+0.512
pragma attribute SERDESIF_075 ment_tsu219 S2_ARADDR[23]->CLK_BASE+0.486
pragma attribute SERDESIF_075 ment_tsu220 S2_ARADDR[24]->CLK_BASE+0.421
pragma attribute SERDESIF_075 ment_tsu221 S2_ARADDR[25]->CLK_BASE+0.764
pragma attribute SERDESIF_075 ment_tsu222 S2_ARADDR[26]->CLK_BASE+0.913
pragma attribute SERDESIF_075 ment_tsu223 S2_ARADDR[27]->CLK_BASE+0.455
pragma attribute SERDESIF_075 ment_tsu224 S2_ARADDR[28]->CLK_BASE+0.996
pragma attribute SERDESIF_075 ment_tsu225 S2_ARADDR[29]->CLK_BASE+0.497
pragma attribute SERDESIF_075 ment_tsu226 S2_ARADDR[2]->CLK_BASE+0.905
pragma attribute SERDESIF_075 ment_tsu227 S2_ARADDR[30]->CLK_BASE+0.309
pragma attribute SERDESIF_075 ment_tsu228 S2_ARADDR[31]->CLK_BASE+0.687
pragma attribute SERDESIF_075 ment_tsu229 S2_ARADDR[3]->CLK_BASE+0.151
pragma attribute SERDESIF_075 ment_tsu230 S2_ARADDR[4]->CLK_BASE+0.344
pragma attribute SERDESIF_075 ment_tsu231 S2_ARADDR[5]->CLK_BASE+0.015
pragma attribute SERDESIF_075 ment_tsu232 S2_ARADDR[6]->CLK_BASE+0.219
pragma attribute SERDESIF_075 ment_tsu233 S2_ARADDR[7]->CLK_BASE+1.025
pragma attribute SERDESIF_075 ment_tsu234 S2_ARADDR[8]->CLK_BASE+0.451
pragma attribute SERDESIF_075 ment_tsu235 S2_ARADDR[9]->CLK_BASE+0.058
pragma attribute SERDESIF_075 ment_tsu236 S2_ARBURST[0]->CLK_BASE+0.517
pragma attribute SERDESIF_075 ment_tsu237 S2_ARBURST[1]->CLK_BASE+0.586
pragma attribute SERDESIF_075 ment_tsu238 S2_ARID[0]->CLK_BASE+0.139
pragma attribute SERDESIF_075 ment_tsu239 S2_ARID[1]->CLK_BASE+0.243
pragma attribute SERDESIF_075 ment_tsu240 S2_ARID[2]->CLK_BASE+0.226
pragma attribute SERDESIF_075 ment_tsu241 S2_ARID[3]->CLK_BASE+0.473
pragma attribute SERDESIF_075 ment_tsu242 S2_ARLEN[0]->CLK_BASE+0.279
pragma attribute SERDESIF_075 ment_tsu243 S2_ARLEN[1]->CLK_BASE+0.540
pragma attribute SERDESIF_075 ment_tsu244 S2_ARLEN[2]->CLK_BASE+0.120
pragma attribute SERDESIF_075 ment_tsu245 S2_ARLEN[3]->CLK_BASE+0.149
pragma attribute SERDESIF_075 ment_tsu246 S2_ARSIZE[0]->CLK_BASE+0.885
pragma attribute SERDESIF_075 ment_tsu247 S2_ARSIZE[1]->CLK_BASE+0.532
pragma attribute SERDESIF_075 ment_tsu248 S2_ARVALID->CLK_BASE+0.392
pragma attribute SERDESIF_075 ment_tsu249 S2_AWADDR_HADDR[0]->CLK_BASE+0.721
pragma attribute SERDESIF_075 ment_tsu250 S2_AWADDR_HADDR[10]->CLK_BASE+0.746
pragma attribute SERDESIF_075 ment_tsu251 S2_AWADDR_HADDR[11]->CLK_BASE+0.568
pragma attribute SERDESIF_075 ment_tsu252 S2_AWADDR_HADDR[12]->CLK_BASE+0.257
pragma attribute SERDESIF_075 ment_tsu253 S2_AWADDR_HADDR[13]->CLK_BASE+0.334
pragma attribute SERDESIF_075 ment_tsu254 S2_AWADDR_HADDR[14]->CLK_BASE+0.446
pragma attribute SERDESIF_075 ment_tsu255 S2_AWADDR_HADDR[15]->CLK_BASE+0.294
pragma attribute SERDESIF_075 ment_tsu256 S2_AWADDR_HADDR[16]->CLK_BASE+0.611
pragma attribute SERDESIF_075 ment_tsu257 S2_AWADDR_HADDR[17]->CLK_BASE+0.435
pragma attribute SERDESIF_075 ment_tsu258 S2_AWADDR_HADDR[18]->CLK_BASE+0.843
pragma attribute SERDESIF_075 ment_tsu259 S2_AWADDR_HADDR[19]->CLK_BASE+0.914
pragma attribute SERDESIF_075 ment_tsu260 S2_AWADDR_HADDR[1]->CLK_BASE+0.464
pragma attribute SERDESIF_075 ment_tsu261 S2_AWADDR_HADDR[20]->CLK_BASE+0.448
pragma attribute SERDESIF_075 ment_tsu262 S2_AWADDR_HADDR[21]->CLK_BASE+0.758
pragma attribute SERDESIF_075 ment_tsu263 S2_AWADDR_HADDR[22]->CLK_BASE+0.672
pragma attribute SERDESIF_075 ment_tsu264 S2_AWADDR_HADDR[23]->CLK_BASE+0.845
pragma attribute SERDESIF_075 ment_tsu265 S2_AWADDR_HADDR[24]->CLK_BASE+0.613
pragma attribute SERDESIF_075 ment_tsu266 S2_AWADDR_HADDR[25]->CLK_BASE+0.650
pragma attribute SERDESIF_075 ment_tsu267 S2_AWADDR_HADDR[26]->CLK_BASE+0.750
pragma attribute SERDESIF_075 ment_tsu268 S2_AWADDR_HADDR[27]->CLK_BASE+0.509
pragma attribute SERDESIF_075 ment_tsu269 S2_AWADDR_HADDR[28]->CLK_BASE+0.672
pragma attribute SERDESIF_075 ment_tsu270 S2_AWADDR_HADDR[29]->CLK_BASE+0.409
pragma attribute SERDESIF_075 ment_tsu271 S2_AWADDR_HADDR[2]->CLK_BASE+0.300
pragma attribute SERDESIF_075 ment_tsu272 S2_AWADDR_HADDR[30]->CLK_BASE+0.933
pragma attribute SERDESIF_075 ment_tsu273 S2_AWADDR_HADDR[31]->CLK_BASE+0.870
pragma attribute SERDESIF_075 ment_tsu274 S2_AWADDR_HADDR[3]->CLK_BASE+0.494
pragma attribute SERDESIF_075 ment_tsu275 S2_AWADDR_HADDR[4]->CLK_BASE+0.640
pragma attribute SERDESIF_075 ment_tsu276 S2_AWADDR_HADDR[5]->CLK_BASE+0.326
pragma attribute SERDESIF_075 ment_tsu277 S2_AWADDR_HADDR[6]->CLK_BASE+0.781
pragma attribute SERDESIF_075 ment_tsu278 S2_AWADDR_HADDR[7]->CLK_BASE+0.341
pragma attribute SERDESIF_075 ment_tsu279 S2_AWADDR_HADDR[8]->CLK_BASE+0.838
pragma attribute SERDESIF_075 ment_tsu280 S2_AWADDR_HADDR[9]->CLK_BASE+0.538
pragma attribute SERDESIF_075 ment_tsu281 S2_AWBURST_HTRANS[0]->CLK_BASE+0.937
pragma attribute SERDESIF_075 ment_tsu282 S2_AWBURST_HTRANS[1]->CLK_BASE+1.035
pragma attribute SERDESIF_075 ment_tsu283 S2_AWID_HSEL[0]->CLK_BASE+1.065
pragma attribute SERDESIF_075 ment_tsu284 S2_AWID_HSEL[1]->CLK_BASE+0.164
pragma attribute SERDESIF_075 ment_tsu285 S2_AWID_HSEL[2]->CLK_BASE+0.109
pragma attribute SERDESIF_075 ment_tsu286 S2_AWID_HSEL[3]->CLK_BASE+-0.015
pragma attribute SERDESIF_075 ment_tsu287 S2_AWLEN_HBURST[0]->CLK_BASE+0.071
pragma attribute SERDESIF_075 ment_tsu288 S2_AWLEN_HBURST[1]->CLK_BASE+-0.029
pragma attribute SERDESIF_075 ment_tsu289 S2_AWLEN_HBURST[2]->CLK_BASE+0.037
pragma attribute SERDESIF_075 ment_tsu290 S2_AWLEN_HBURST[3]->CLK_BASE+0.425
pragma attribute SERDESIF_075 ment_tsu291 S2_AWSIZE_HSIZE[0]->CLK_BASE+0.939
pragma attribute SERDESIF_075 ment_tsu292 S2_AWSIZE_HSIZE[1]->CLK_BASE+0.740
pragma attribute SERDESIF_075 ment_tsu293 S2_AWVALID_HWRITE->CLK_BASE+0.798
pragma attribute SERDESIF_075 ment_tsu294 S2_BREADY_HREADY->CLK_BASE+0.972
pragma attribute SERDESIF_075 ment_tsu295 S2_RREADY->CLK_BASE+0.850
pragma attribute SERDESIF_075 ment_tsu296 S2_WDATA_HWDATA[0]->CLK_BASE+0.007
pragma attribute SERDESIF_075 ment_tsu297 S2_WDATA_HWDATA[10]->CLK_BASE+0.147
pragma attribute SERDESIF_075 ment_tsu298 S2_WDATA_HWDATA[11]->CLK_BASE+0.088
pragma attribute SERDESIF_075 ment_tsu299 S2_WDATA_HWDATA[12]->CLK_BASE+0.187
pragma attribute SERDESIF_075 ment_tsu300 S2_WDATA_HWDATA[13]->CLK_BASE+0.242
pragma attribute SERDESIF_075 ment_tsu301 S2_WDATA_HWDATA[14]->CLK_BASE+0.179
pragma attribute SERDESIF_075 ment_tsu302 S2_WDATA_HWDATA[15]->CLK_BASE+0.120
pragma attribute SERDESIF_075 ment_tsu303 S2_WDATA_HWDATA[16]->CLK_BASE+0.108
pragma attribute SERDESIF_075 ment_tsu304 S2_WDATA_HWDATA[17]->CLK_BASE+0.173
pragma attribute SERDESIF_075 ment_tsu305 S2_WDATA_HWDATA[18]->CLK_BASE+0.427
pragma attribute SERDESIF_075 ment_tsu306 S2_WDATA_HWDATA[19]->CLK_BASE+0.236
pragma attribute SERDESIF_075 ment_tsu307 S2_WDATA_HWDATA[1]->CLK_BASE+0.051
pragma attribute SERDESIF_075 ment_tsu308 S2_WDATA_HWDATA[20]->CLK_BASE+0.281
pragma attribute SERDESIF_075 ment_tsu309 S2_WDATA_HWDATA[21]->CLK_BASE+-0.045
pragma attribute SERDESIF_075 ment_tsu310 S2_WDATA_HWDATA[22]->CLK_BASE+0.144
pragma attribute SERDESIF_075 ment_tsu311 S2_WDATA_HWDATA[23]->CLK_BASE+0.163
pragma attribute SERDESIF_075 ment_tsu312 S2_WDATA_HWDATA[24]->CLK_BASE+0.324
pragma attribute SERDESIF_075 ment_tsu313 S2_WDATA_HWDATA[25]->CLK_BASE+0.307
pragma attribute SERDESIF_075 ment_tsu314 S2_WDATA_HWDATA[26]->CLK_BASE+0.169
pragma attribute SERDESIF_075 ment_tsu315 S2_WDATA_HWDATA[27]->CLK_BASE+0.185
pragma attribute SERDESIF_075 ment_tsu316 S2_WDATA_HWDATA[28]->CLK_BASE+0.436
pragma attribute SERDESIF_075 ment_tsu317 S2_WDATA_HWDATA[29]->CLK_BASE+0.353
pragma attribute SERDESIF_075 ment_tsu318 S2_WDATA_HWDATA[2]->CLK_BASE+0.136
pragma attribute SERDESIF_075 ment_tsu319 S2_WDATA_HWDATA[30]->CLK_BASE+0.152
pragma attribute SERDESIF_075 ment_tsu320 S2_WDATA_HWDATA[31]->CLK_BASE+0.288
pragma attribute SERDESIF_075 ment_tsu321 S2_WDATA_HWDATA[32]->CLK_BASE+0.190
pragma attribute SERDESIF_075 ment_tsu322 S2_WDATA_HWDATA[33]->CLK_BASE+0.555
pragma attribute SERDESIF_075 ment_tsu323 S2_WDATA_HWDATA[34]->CLK_BASE+0.466
pragma attribute SERDESIF_075 ment_tsu324 S2_WDATA_HWDATA[35]->CLK_BASE+0.424
pragma attribute SERDESIF_075 ment_tsu325 S2_WDATA_HWDATA[36]->CLK_BASE+0.212
pragma attribute SERDESIF_075 ment_tsu326 S2_WDATA_HWDATA[37]->CLK_BASE+0.026
pragma attribute SERDESIF_075 ment_tsu327 S2_WDATA_HWDATA[38]->CLK_BASE+0.004
pragma attribute SERDESIF_075 ment_tsu328 S2_WDATA_HWDATA[39]->CLK_BASE+-0.032
pragma attribute SERDESIF_075 ment_tsu329 S2_WDATA_HWDATA[3]->CLK_BASE+0.044
pragma attribute SERDESIF_075 ment_tsu330 S2_WDATA_HWDATA[40]->CLK_BASE+-0.023
pragma attribute SERDESIF_075 ment_tsu331 S2_WDATA_HWDATA[41]->CLK_BASE+-0.063
pragma attribute SERDESIF_075 ment_tsu332 S2_WDATA_HWDATA[42]->CLK_BASE+0.447
pragma attribute SERDESIF_075 ment_tsu333 S2_WDATA_HWDATA[43]->CLK_BASE+0.703
pragma attribute SERDESIF_075 ment_tsu334 S2_WDATA_HWDATA[44]->CLK_BASE+-0.033
pragma attribute SERDESIF_075 ment_tsu335 S2_WDATA_HWDATA[45]->CLK_BASE+0.037
pragma attribute SERDESIF_075 ment_tsu336 S2_WDATA_HWDATA[46]->CLK_BASE+0.295
pragma attribute SERDESIF_075 ment_tsu337 S2_WDATA_HWDATA[47]->CLK_BASE+-0.039
pragma attribute SERDESIF_075 ment_tsu338 S2_WDATA_HWDATA[48]->CLK_BASE+0.505
pragma attribute SERDESIF_075 ment_tsu339 S2_WDATA_HWDATA[49]->CLK_BASE+0.176
pragma attribute SERDESIF_075 ment_tsu340 S2_WDATA_HWDATA[4]->CLK_BASE+0.380
pragma attribute SERDESIF_075 ment_tsu341 S2_WDATA_HWDATA[50]->CLK_BASE+0.269
pragma attribute SERDESIF_075 ment_tsu342 S2_WDATA_HWDATA[51]->CLK_BASE+0.110
pragma attribute SERDESIF_075 ment_tsu343 S2_WDATA_HWDATA[52]->CLK_BASE+0.046
pragma attribute SERDESIF_075 ment_tsu344 S2_WDATA_HWDATA[53]->CLK_BASE+-0.054
pragma attribute SERDESIF_075 ment_tsu345 S2_WDATA_HWDATA[54]->CLK_BASE+0.045
pragma attribute SERDESIF_075 ment_tsu346 S2_WDATA_HWDATA[55]->CLK_BASE+-0.163
pragma attribute SERDESIF_075 ment_tsu347 S2_WDATA_HWDATA[56]->CLK_BASE+0.423
pragma attribute SERDESIF_075 ment_tsu348 S2_WDATA_HWDATA[57]->CLK_BASE+0.370
pragma attribute SERDESIF_075 ment_tsu349 S2_WDATA_HWDATA[58]->CLK_BASE+0.004
pragma attribute SERDESIF_075 ment_tsu350 S2_WDATA_HWDATA[59]->CLK_BASE+-0.182
pragma attribute SERDESIF_075 ment_tsu351 S2_WDATA_HWDATA[5]->CLK_BASE+0.432
pragma attribute SERDESIF_075 ment_tsu352 S2_WDATA_HWDATA[60]->CLK_BASE+0.046
pragma attribute SERDESIF_075 ment_tsu353 S2_WDATA_HWDATA[61]->CLK_BASE+-0.133
pragma attribute SERDESIF_075 ment_tsu354 S2_WDATA_HWDATA[62]->CLK_BASE+0.428
pragma attribute SERDESIF_075 ment_tsu355 S2_WDATA_HWDATA[63]->CLK_BASE+0.148
pragma attribute SERDESIF_075 ment_tsu356 S2_WDATA_HWDATA[6]->CLK_BASE+0.137
pragma attribute SERDESIF_075 ment_tsu357 S2_WDATA_HWDATA[7]->CLK_BASE+0.407
pragma attribute SERDESIF_075 ment_tsu358 S2_WDATA_HWDATA[8]->CLK_BASE+0.669
pragma attribute SERDESIF_075 ment_tsu359 S2_WDATA_HWDATA[9]->CLK_BASE+0.093
pragma attribute SERDESIF_075 ment_tsu360 S2_WLAST->CLK_BASE+0.265
pragma attribute SERDESIF_075 ment_tsu361 S2_WSTRB[0]->CLK_BASE+0.685
pragma attribute SERDESIF_075 ment_tsu362 S2_WSTRB[1]->CLK_BASE+0.313
pragma attribute SERDESIF_075 ment_tsu363 S2_WSTRB[2]->CLK_BASE+0.535
pragma attribute SERDESIF_075 ment_tsu364 S2_WSTRB[3]->CLK_BASE+0.323
pragma attribute SERDESIF_075 ment_tsu365 S2_WSTRB[4]->CLK_BASE+0.083
pragma attribute SERDESIF_075 ment_tsu366 S2_WSTRB[5]->CLK_BASE+0.671
pragma attribute SERDESIF_075 ment_tsu367 S2_WSTRB[6]->CLK_BASE+0.424
pragma attribute SERDESIF_075 ment_tsu368 S2_WSTRB[7]->CLK_BASE+0.391
pragma attribute SERDESIF_075 ment_tsu369 S2_WVALID->CLK_BASE+0.437
pragma attribute SERDESIF_075 ment_tsu370 S_ARADDR[0]->CLK_BASE+0.852
pragma attribute SERDESIF_075 ment_tsu371 S_ARADDR[10]->CLK_BASE+1.011
pragma attribute SERDESIF_075 ment_tsu372 S_ARADDR[11]->CLK_BASE+0.989
pragma attribute SERDESIF_075 ment_tsu373 S_ARADDR[12]->CLK_BASE+0.622
pragma attribute SERDESIF_075 ment_tsu374 S_ARADDR[13]->CLK_BASE+0.694
pragma attribute SERDESIF_075 ment_tsu375 S_ARADDR[14]->CLK_BASE+0.938
pragma attribute SERDESIF_075 ment_tsu376 S_ARADDR[15]->CLK_BASE+0.545
pragma attribute SERDESIF_075 ment_tsu377 S_ARADDR[16]->CLK_BASE+0.513
pragma attribute SERDESIF_075 ment_tsu378 S_ARADDR[17]->CLK_BASE+0.871
pragma attribute SERDESIF_075 ment_tsu379 S_ARADDR[18]->CLK_BASE+1.032
pragma attribute SERDESIF_075 ment_tsu380 S_ARADDR[19]->CLK_BASE+0.883
pragma attribute SERDESIF_075 ment_tsu381 S_ARADDR[1]->CLK_BASE+0.420
pragma attribute SERDESIF_075 ment_tsu382 S_ARADDR[20]->CLK_BASE+0.873
pragma attribute SERDESIF_075 ment_tsu383 S_ARADDR[21]->CLK_BASE+0.757
pragma attribute SERDESIF_075 ment_tsu384 S_ARADDR[22]->CLK_BASE+0.761
pragma attribute SERDESIF_075 ment_tsu385 S_ARADDR[23]->CLK_BASE+0.942
pragma attribute SERDESIF_075 ment_tsu386 S_ARADDR[24]->CLK_BASE+0.556
pragma attribute SERDESIF_075 ment_tsu387 S_ARADDR[25]->CLK_BASE+0.594
pragma attribute SERDESIF_075 ment_tsu388 S_ARADDR[26]->CLK_BASE+0.599
pragma attribute SERDESIF_075 ment_tsu389 S_ARADDR[27]->CLK_BASE+0.923
pragma attribute SERDESIF_075 ment_tsu390 S_ARADDR[28]->CLK_BASE+0.588
pragma attribute SERDESIF_075 ment_tsu391 S_ARADDR[29]->CLK_BASE+0.713
pragma attribute SERDESIF_075 ment_tsu392 S_ARADDR[2]->CLK_BASE+0.736
pragma attribute SERDESIF_075 ment_tsu393 S_ARADDR[30]->CLK_BASE+0.680
pragma attribute SERDESIF_075 ment_tsu394 S_ARADDR[31]->CLK_BASE+0.659
pragma attribute SERDESIF_075 ment_tsu395 S_ARADDR[3]->CLK_BASE+1.077
pragma attribute SERDESIF_075 ment_tsu396 S_ARADDR[4]->CLK_BASE+0.514
pragma attribute SERDESIF_075 ment_tsu397 S_ARADDR[5]->CLK_BASE+0.678
pragma attribute SERDESIF_075 ment_tsu398 S_ARADDR[6]->CLK_BASE+1.054
pragma attribute SERDESIF_075 ment_tsu399 S_ARADDR[7]->CLK_BASE+0.686
pragma attribute SERDESIF_075 ment_tsu400 S_ARADDR[8]->CLK_BASE+0.971
pragma attribute SERDESIF_075 ment_tsu401 S_ARADDR[9]->CLK_BASE+0.791
pragma attribute SERDESIF_075 ment_tsu402 S_ARBURST[0]->CLK_BASE+0.564
pragma attribute SERDESIF_075 ment_tsu403 S_ARBURST[1]->CLK_BASE+0.491
pragma attribute SERDESIF_075 ment_tsu404 S_ARID[0]->CLK_BASE+0.656
pragma attribute SERDESIF_075 ment_tsu405 S_ARID[1]->CLK_BASE+0.647
pragma attribute SERDESIF_075 ment_tsu406 S_ARID[2]->CLK_BASE+0.708
pragma attribute SERDESIF_075 ment_tsu407 S_ARID[3]->CLK_BASE+0.638
pragma attribute SERDESIF_075 ment_tsu408 S_ARLEN[0]->CLK_BASE+0.569
pragma attribute SERDESIF_075 ment_tsu409 S_ARLEN[1]->CLK_BASE+0.659
pragma attribute SERDESIF_075 ment_tsu410 S_ARLEN[2]->CLK_BASE+0.607
pragma attribute SERDESIF_075 ment_tsu411 S_ARLEN[3]->CLK_BASE+0.511
pragma attribute SERDESIF_075 ment_tsu412 S_ARSIZE[0]->CLK_BASE+0.618
pragma attribute SERDESIF_075 ment_tsu413 S_ARSIZE[1]->CLK_BASE+0.896
pragma attribute SERDESIF_075 ment_tsu414 S_ARVALID->CLK_BASE+0.664
pragma attribute SERDESIF_075 ment_tsu415 S_AWADDR_HADDR[0]->CLK_BASE+0.622
pragma attribute SERDESIF_075 ment_tsu416 S_AWADDR_HADDR[10]->CLK_BASE+0.797
pragma attribute SERDESIF_075 ment_tsu417 S_AWADDR_HADDR[11]->CLK_BASE+0.933
pragma attribute SERDESIF_075 ment_tsu418 S_AWADDR_HADDR[12]->CLK_BASE+0.739
pragma attribute SERDESIF_075 ment_tsu419 S_AWADDR_HADDR[13]->CLK_BASE+0.878
pragma attribute SERDESIF_075 ment_tsu420 S_AWADDR_HADDR[14]->CLK_BASE+0.821
pragma attribute SERDESIF_075 ment_tsu421 S_AWADDR_HADDR[15]->CLK_BASE+0.614
pragma attribute SERDESIF_075 ment_tsu422 S_AWADDR_HADDR[16]->CLK_BASE+0.704
pragma attribute SERDESIF_075 ment_tsu423 S_AWADDR_HADDR[17]->CLK_BASE+0.839
pragma attribute SERDESIF_075 ment_tsu424 S_AWADDR_HADDR[18]->CLK_BASE+1.037
pragma attribute SERDESIF_075 ment_tsu425 S_AWADDR_HADDR[19]->CLK_BASE+0.748
pragma attribute SERDESIF_075 ment_tsu426 S_AWADDR_HADDR[1]->CLK_BASE+0.677
pragma attribute SERDESIF_075 ment_tsu427 S_AWADDR_HADDR[20]->CLK_BASE+0.727
pragma attribute SERDESIF_075 ment_tsu428 S_AWADDR_HADDR[21]->CLK_BASE+0.819
pragma attribute SERDESIF_075 ment_tsu429 S_AWADDR_HADDR[22]->CLK_BASE+0.886
pragma attribute SERDESIF_075 ment_tsu430 S_AWADDR_HADDR[23]->CLK_BASE+0.760
pragma attribute SERDESIF_075 ment_tsu431 S_AWADDR_HADDR[24]->CLK_BASE+0.630
pragma attribute SERDESIF_075 ment_tsu432 S_AWADDR_HADDR[25]->CLK_BASE+0.972
pragma attribute SERDESIF_075 ment_tsu433 S_AWADDR_HADDR[26]->CLK_BASE+0.513
pragma attribute SERDESIF_075 ment_tsu434 S_AWADDR_HADDR[27]->CLK_BASE+0.890
pragma attribute SERDESIF_075 ment_tsu435 S_AWADDR_HADDR[28]->CLK_BASE+0.670
pragma attribute SERDESIF_075 ment_tsu436 S_AWADDR_HADDR[29]->CLK_BASE+0.900
pragma attribute SERDESIF_075 ment_tsu437 S_AWADDR_HADDR[2]->CLK_BASE+0.612
pragma attribute SERDESIF_075 ment_tsu438 S_AWADDR_HADDR[30]->CLK_BASE+0.884
pragma attribute SERDESIF_075 ment_tsu439 S_AWADDR_HADDR[31]->CLK_BASE+0.751
pragma attribute SERDESIF_075 ment_tsu440 S_AWADDR_HADDR[3]->CLK_BASE+0.924
pragma attribute SERDESIF_075 ment_tsu441 S_AWADDR_HADDR[4]->CLK_BASE+0.584
pragma attribute SERDESIF_075 ment_tsu442 S_AWADDR_HADDR[5]->CLK_BASE+0.479
pragma attribute SERDESIF_075 ment_tsu443 S_AWADDR_HADDR[6]->CLK_BASE+0.650
pragma attribute SERDESIF_075 ment_tsu444 S_AWADDR_HADDR[7]->CLK_BASE+0.937
pragma attribute SERDESIF_075 ment_tsu445 S_AWADDR_HADDR[8]->CLK_BASE+0.454
pragma attribute SERDESIF_075 ment_tsu446 S_AWADDR_HADDR[9]->CLK_BASE+0.665
pragma attribute SERDESIF_075 ment_tsu447 S_AWBURST_HTRANS[0]->CLK_BASE+0.862
pragma attribute SERDESIF_075 ment_tsu448 S_AWBURST_HTRANS[1]->CLK_BASE+0.881
pragma attribute SERDESIF_075 ment_tsu449 S_AWID_HSEL[0]->CLK_BASE+0.793
pragma attribute SERDESIF_075 ment_tsu450 S_AWID_HSEL[1]->CLK_BASE+0.460
pragma attribute SERDESIF_075 ment_tsu451 S_AWID_HSEL[2]->CLK_BASE+0.422
pragma attribute SERDESIF_075 ment_tsu452 S_AWID_HSEL[3]->CLK_BASE+0.245
pragma attribute SERDESIF_075 ment_tsu453 S_AWLEN_HBURST[0]->CLK_BASE+0.530
pragma attribute SERDESIF_075 ment_tsu454 S_AWLEN_HBURST[1]->CLK_BASE+0.207
pragma attribute SERDESIF_075 ment_tsu455 S_AWLEN_HBURST[2]->CLK_BASE+0.582
pragma attribute SERDESIF_075 ment_tsu456 S_AWLEN_HBURST[3]->CLK_BASE+0.649
pragma attribute SERDESIF_075 ment_tsu457 S_AWSIZE_HSIZE[0]->CLK_BASE+0.996
pragma attribute SERDESIF_075 ment_tsu458 S_AWSIZE_HSIZE[1]->CLK_BASE+0.963
pragma attribute SERDESIF_075 ment_tsu459 S_AWVALID_HWRITE->CLK_BASE+0.783
pragma attribute SERDESIF_075 ment_tsu460 S_BREADY_HREADY->CLK_BASE+1.046
pragma attribute SERDESIF_075 ment_tsu461 S_RREADY->CLK_BASE+0.878
pragma attribute SERDESIF_075 ment_tsu462 S_WDATA_HWDATA[0]->CLK_BASE+0.548
pragma attribute SERDESIF_075 ment_tsu463 S_WDATA_HWDATA[10]->CLK_BASE+0.273
pragma attribute SERDESIF_075 ment_tsu464 S_WDATA_HWDATA[11]->CLK_BASE+0.544
pragma attribute SERDESIF_075 ment_tsu465 S_WDATA_HWDATA[12]->CLK_BASE+0.351
pragma attribute SERDESIF_075 ment_tsu466 S_WDATA_HWDATA[13]->CLK_BASE+0.607
pragma attribute SERDESIF_075 ment_tsu467 S_WDATA_HWDATA[14]->CLK_BASE+0.284
pragma attribute SERDESIF_075 ment_tsu468 S_WDATA_HWDATA[15]->CLK_BASE+0.328
pragma attribute SERDESIF_075 ment_tsu469 S_WDATA_HWDATA[16]->CLK_BASE+0.379
pragma attribute SERDESIF_075 ment_tsu470 S_WDATA_HWDATA[17]->CLK_BASE+0.668
pragma attribute SERDESIF_075 ment_tsu471 S_WDATA_HWDATA[18]->CLK_BASE+0.496
pragma attribute SERDESIF_075 ment_tsu472 S_WDATA_HWDATA[19]->CLK_BASE+0.333
pragma attribute SERDESIF_075 ment_tsu473 S_WDATA_HWDATA[1]->CLK_BASE+0.646
pragma attribute SERDESIF_075 ment_tsu474 S_WDATA_HWDATA[20]->CLK_BASE+0.381
pragma attribute SERDESIF_075 ment_tsu475 S_WDATA_HWDATA[21]->CLK_BASE+0.462
pragma attribute SERDESIF_075 ment_tsu476 S_WDATA_HWDATA[22]->CLK_BASE+0.320
pragma attribute SERDESIF_075 ment_tsu477 S_WDATA_HWDATA[23]->CLK_BASE+0.621
pragma attribute SERDESIF_075 ment_tsu478 S_WDATA_HWDATA[24]->CLK_BASE+0.258
pragma attribute SERDESIF_075 ment_tsu479 S_WDATA_HWDATA[25]->CLK_BASE+0.380
pragma attribute SERDESIF_075 ment_tsu480 S_WDATA_HWDATA[26]->CLK_BASE+0.529
pragma attribute SERDESIF_075 ment_tsu481 S_WDATA_HWDATA[27]->CLK_BASE+0.659
pragma attribute SERDESIF_075 ment_tsu482 S_WDATA_HWDATA[28]->CLK_BASE+0.334
pragma attribute SERDESIF_075 ment_tsu483 S_WDATA_HWDATA[29]->CLK_BASE+0.546
pragma attribute SERDESIF_075 ment_tsu484 S_WDATA_HWDATA[2]->CLK_BASE+0.241
pragma attribute SERDESIF_075 ment_tsu485 S_WDATA_HWDATA[30]->CLK_BASE+0.245
pragma attribute SERDESIF_075 ment_tsu486 S_WDATA_HWDATA[31]->CLK_BASE+0.684
pragma attribute SERDESIF_075 ment_tsu487 S_WDATA_HWDATA[32]->CLK_BASE+0.658
pragma attribute SERDESIF_075 ment_tsu488 S_WDATA_HWDATA[33]->CLK_BASE+0.712
pragma attribute SERDESIF_075 ment_tsu489 S_WDATA_HWDATA[34]->CLK_BASE+0.726
pragma attribute SERDESIF_075 ment_tsu490 S_WDATA_HWDATA[35]->CLK_BASE+0.756
pragma attribute SERDESIF_075 ment_tsu491 S_WDATA_HWDATA[36]->CLK_BASE+0.301
pragma attribute SERDESIF_075 ment_tsu492 S_WDATA_HWDATA[37]->CLK_BASE+0.562
pragma attribute SERDESIF_075 ment_tsu493 S_WDATA_HWDATA[38]->CLK_BASE+0.715
pragma attribute SERDESIF_075 ment_tsu494 S_WDATA_HWDATA[39]->CLK_BASE+0.520
pragma attribute SERDESIF_075 ment_tsu495 S_WDATA_HWDATA[3]->CLK_BASE+0.288
pragma attribute SERDESIF_075 ment_tsu496 S_WDATA_HWDATA[40]->CLK_BASE+0.297
pragma attribute SERDESIF_075 ment_tsu497 S_WDATA_HWDATA[41]->CLK_BASE+0.524
pragma attribute SERDESIF_075 ment_tsu498 S_WDATA_HWDATA[42]->CLK_BASE+0.723
pragma attribute SERDESIF_075 ment_tsu499 S_WDATA_HWDATA[43]->CLK_BASE+0.715
pragma attribute SERDESIF_075 ment_tsu500 S_WDATA_HWDATA[44]->CLK_BASE+0.353
pragma attribute SERDESIF_075 ment_tsu501 S_WDATA_HWDATA[45]->CLK_BASE+0.349
pragma attribute SERDESIF_075 ment_tsu502 S_WDATA_HWDATA[46]->CLK_BASE+0.783
pragma attribute SERDESIF_075 ment_tsu503 S_WDATA_HWDATA[47]->CLK_BASE+0.467
pragma attribute SERDESIF_075 ment_tsu504 S_WDATA_HWDATA[48]->CLK_BASE+0.519
pragma attribute SERDESIF_075 ment_tsu505 S_WDATA_HWDATA[49]->CLK_BASE+0.336
pragma attribute SERDESIF_075 ment_tsu506 S_WDATA_HWDATA[4]->CLK_BASE+0.231
pragma attribute SERDESIF_075 ment_tsu507 S_WDATA_HWDATA[50]->CLK_BASE+0.340
pragma attribute SERDESIF_075 ment_tsu508 S_WDATA_HWDATA[51]->CLK_BASE+0.747
pragma attribute SERDESIF_075 ment_tsu509 S_WDATA_HWDATA[52]->CLK_BASE+0.578
pragma attribute SERDESIF_075 ment_tsu510 S_WDATA_HWDATA[53]->CLK_BASE+0.664
pragma attribute SERDESIF_075 ment_tsu511 S_WDATA_HWDATA[54]->CLK_BASE+0.690
pragma attribute SERDESIF_075 ment_tsu512 S_WDATA_HWDATA[55]->CLK_BASE+0.567
pragma attribute SERDESIF_075 ment_tsu513 S_WDATA_HWDATA[56]->CLK_BASE+0.752
pragma attribute SERDESIF_075 ment_tsu514 S_WDATA_HWDATA[57]->CLK_BASE+0.560
pragma attribute SERDESIF_075 ment_tsu515 S_WDATA_HWDATA[58]->CLK_BASE+0.541
pragma attribute SERDESIF_075 ment_tsu516 S_WDATA_HWDATA[59]->CLK_BASE+0.487
pragma attribute SERDESIF_075 ment_tsu517 S_WDATA_HWDATA[5]->CLK_BASE+0.253
pragma attribute SERDESIF_075 ment_tsu518 S_WDATA_HWDATA[60]->CLK_BASE+0.580
pragma attribute SERDESIF_075 ment_tsu519 S_WDATA_HWDATA[61]->CLK_BASE+0.552
pragma attribute SERDESIF_075 ment_tsu520 S_WDATA_HWDATA[62]->CLK_BASE+0.291
pragma attribute SERDESIF_075 ment_tsu521 S_WDATA_HWDATA[63]->CLK_BASE+0.530
pragma attribute SERDESIF_075 ment_tsu522 S_WDATA_HWDATA[6]->CLK_BASE+0.631
pragma attribute SERDESIF_075 ment_tsu523 S_WDATA_HWDATA[7]->CLK_BASE+0.726
pragma attribute SERDESIF_075 ment_tsu524 S_WDATA_HWDATA[8]->CLK_BASE+0.303
pragma attribute SERDESIF_075 ment_tsu525 S_WDATA_HWDATA[9]->CLK_BASE+0.320
pragma attribute SERDESIF_075 ment_tsu526 S_WLAST->CLK_BASE+0.467
pragma attribute SERDESIF_075 ment_tsu527 S_WSTRB[0]->CLK_BASE+0.711
pragma attribute SERDESIF_075 ment_tsu528 S_WSTRB[1]->CLK_BASE+0.827
pragma attribute SERDESIF_075 ment_tsu529 S_WSTRB[2]->CLK_BASE+0.955
pragma attribute SERDESIF_075 ment_tsu530 S_WSTRB[3]->CLK_BASE+0.862
pragma attribute SERDESIF_075 ment_tsu531 S_WSTRB[4]->CLK_BASE+0.537
pragma attribute SERDESIF_075 ment_tsu532 S_WSTRB[5]->CLK_BASE+0.910
pragma attribute SERDESIF_075 ment_tsu533 S_WSTRB[6]->CLK_BASE+0.403
pragma attribute SERDESIF_075 ment_tsu534 S_WSTRB[7]->CLK_BASE+0.633
pragma attribute SERDESIF_075 ment_tsu535 S_WVALID->CLK_BASE+0.703
pragma attribute SERDESIF_075 ment_tco0 APB_CLK->APB_PRDATA[0]+4.934
pragma attribute SERDESIF_075 ment_tco1 APB_CLK->APB_PRDATA[10]+5.024
pragma attribute SERDESIF_075 ment_tco2 APB_CLK->APB_PRDATA[11]+5.105
pragma attribute SERDESIF_075 ment_tco3 APB_CLK->APB_PRDATA[12]+5.156
pragma attribute SERDESIF_075 ment_tco4 APB_CLK->APB_PRDATA[13]+5.196
pragma attribute SERDESIF_075 ment_tco5 APB_CLK->APB_PRDATA[14]+5.014
pragma attribute SERDESIF_075 ment_tco6 APB_CLK->APB_PRDATA[15]+5.106
pragma attribute SERDESIF_075 ment_tco7 APB_CLK->APB_PRDATA[16]+5.048
pragma attribute SERDESIF_075 ment_tco8 APB_CLK->APB_PRDATA[17]+5.201
pragma attribute SERDESIF_075 ment_tco9 APB_CLK->APB_PRDATA[18]+5.007
pragma attribute SERDESIF_075 ment_tco10 APB_CLK->APB_PRDATA[19]+5.160
pragma attribute SERDESIF_075 ment_tco11 APB_CLK->APB_PRDATA[1]+4.896
pragma attribute SERDESIF_075 ment_tco12 APB_CLK->APB_PRDATA[20]+5.049
pragma attribute SERDESIF_075 ment_tco13 APB_CLK->APB_PRDATA[21]+5.157
pragma attribute SERDESIF_075 ment_tco14 APB_CLK->APB_PRDATA[22]+5.029
pragma attribute SERDESIF_075 ment_tco15 APB_CLK->APB_PRDATA[23]+5.161
pragma attribute SERDESIF_075 ment_tco16 APB_CLK->APB_PRDATA[24]+5.230
pragma attribute SERDESIF_075 ment_tco17 APB_CLK->APB_PRDATA[25]+5.348
pragma attribute SERDESIF_075 ment_tco18 APB_CLK->APB_PRDATA[26]+5.076
pragma attribute SERDESIF_075 ment_tco19 APB_CLK->APB_PRDATA[27]+5.125
pragma attribute SERDESIF_075 ment_tco20 APB_CLK->APB_PRDATA[28]+5.217
pragma attribute SERDESIF_075 ment_tco21 APB_CLK->APB_PRDATA[29]+5.235
pragma attribute SERDESIF_075 ment_tco22 APB_CLK->APB_PRDATA[2]+5.014
pragma attribute SERDESIF_075 ment_tco23 APB_CLK->APB_PRDATA[30]+4.986
pragma attribute SERDESIF_075 ment_tco24 APB_CLK->APB_PRDATA[31]+5.038
pragma attribute SERDESIF_075 ment_tco25 APB_CLK->APB_PRDATA[3]+4.838
pragma attribute SERDESIF_075 ment_tco26 APB_CLK->APB_PRDATA[4]+4.918
pragma attribute SERDESIF_075 ment_tco27 APB_CLK->APB_PRDATA[5]+4.908
pragma attribute SERDESIF_075 ment_tco28 APB_CLK->APB_PRDATA[6]+4.814
pragma attribute SERDESIF_075 ment_tco29 APB_CLK->APB_PRDATA[7]+4.869
pragma attribute SERDESIF_075 ment_tco30 APB_CLK->APB_PRDATA[8]+5.255
pragma attribute SERDESIF_075 ment_tco31 APB_CLK->APB_PRDATA[9]+5.129
pragma attribute SERDESIF_075 ment_tco32 APB_CLK->APB_PREADY+4.732
pragma attribute SERDESIF_075 ment_tco33 APB_CLK->APB_PSLVERR+4.957
pragma attribute SERDESIF_075 ment_tco34 APB_CLK->PCIE2_SYSTEM_INT+3.792
pragma attribute SERDESIF_075 ment_tco35 APB_CLK->PCIE_SYSTEM_INT+4.040
pragma attribute SERDESIF_075 ment_tco36 APB_CLK->PLL_LOCKLOST_INT+3.655
pragma attribute SERDESIF_075 ment_tco37 APB_CLK->PLL_LOCK_INT+3.873
pragma attribute SERDESIF_075 ment_tco38 CLK_BASE->M2_ARADDR[0]+3.154
pragma attribute SERDESIF_075 ment_tco39 CLK_BASE->M2_ARADDR[10]+3.207
pragma attribute SERDESIF_075 ment_tco40 CLK_BASE->M2_ARADDR[11]+3.120
pragma attribute SERDESIF_075 ment_tco41 CLK_BASE->M2_ARADDR[12]+3.218
pragma attribute SERDESIF_075 ment_tco42 CLK_BASE->M2_ARADDR[13]+3.227
pragma attribute SERDESIF_075 ment_tco43 CLK_BASE->M2_ARADDR[14]+3.268
pragma attribute SERDESIF_075 ment_tco44 CLK_BASE->M2_ARADDR[15]+3.253
pragma attribute SERDESIF_075 ment_tco45 CLK_BASE->M2_ARADDR[16]+3.215
pragma attribute SERDESIF_075 ment_tco46 CLK_BASE->M2_ARADDR[17]+3.229
pragma attribute SERDESIF_075 ment_tco47 CLK_BASE->M2_ARADDR[18]+3.184
pragma attribute SERDESIF_075 ment_tco48 CLK_BASE->M2_ARADDR[19]+3.181
pragma attribute SERDESIF_075 ment_tco49 CLK_BASE->M2_ARADDR[1]+3.133
pragma attribute SERDESIF_075 ment_tco50 CLK_BASE->M2_ARADDR[20]+3.125
pragma attribute SERDESIF_075 ment_tco51 CLK_BASE->M2_ARADDR[21]+3.251
pragma attribute SERDESIF_075 ment_tco52 CLK_BASE->M2_ARADDR[22]+3.190
pragma attribute SERDESIF_075 ment_tco53 CLK_BASE->M2_ARADDR[23]+3.229
pragma attribute SERDESIF_075 ment_tco54 CLK_BASE->M2_ARADDR[24]+3.238
pragma attribute SERDESIF_075 ment_tco55 CLK_BASE->M2_ARADDR[25]+3.071
pragma attribute SERDESIF_075 ment_tco56 CLK_BASE->M2_ARADDR[26]+3.105
pragma attribute SERDESIF_075 ment_tco57 CLK_BASE->M2_ARADDR[27]+3.206
pragma attribute SERDESIF_075 ment_tco58 CLK_BASE->M2_ARADDR[28]+3.191
pragma attribute SERDESIF_075 ment_tco59 CLK_BASE->M2_ARADDR[29]+3.127
pragma attribute SERDESIF_075 ment_tco60 CLK_BASE->M2_ARADDR[2]+3.180
pragma attribute SERDESIF_075 ment_tco61 CLK_BASE->M2_ARADDR[30]+3.080
pragma attribute SERDESIF_075 ment_tco62 CLK_BASE->M2_ARADDR[31]+3.207
pragma attribute SERDESIF_075 ment_tco63 CLK_BASE->M2_ARADDR[3]+3.130
pragma attribute SERDESIF_075 ment_tco64 CLK_BASE->M2_ARADDR[4]+3.135
pragma attribute SERDESIF_075 ment_tco65 CLK_BASE->M2_ARADDR[5]+3.116
pragma attribute SERDESIF_075 ment_tco66 CLK_BASE->M2_ARADDR[6]+3.218
pragma attribute SERDESIF_075 ment_tco67 CLK_BASE->M2_ARADDR[7]+3.150
pragma attribute SERDESIF_075 ment_tco68 CLK_BASE->M2_ARADDR[8]+3.163
pragma attribute SERDESIF_075 ment_tco69 CLK_BASE->M2_ARADDR[9]+3.256
pragma attribute SERDESIF_075 ment_tco70 CLK_BASE->M2_ARBURST[0]+3.128
pragma attribute SERDESIF_075 ment_tco71 CLK_BASE->M2_ARID[0]+3.117
pragma attribute SERDESIF_075 ment_tco72 CLK_BASE->M2_ARID[1]+3.094
pragma attribute SERDESIF_075 ment_tco73 CLK_BASE->M2_ARLEN[0]+3.156
pragma attribute SERDESIF_075 ment_tco74 CLK_BASE->M2_ARLEN[1]+3.137
pragma attribute SERDESIF_075 ment_tco75 CLK_BASE->M2_ARLEN[2]+3.086
pragma attribute SERDESIF_075 ment_tco76 CLK_BASE->M2_ARLEN[3]+3.112
pragma attribute SERDESIF_075 ment_tco77 CLK_BASE->M2_ARSIZE[0]+3.176
pragma attribute SERDESIF_075 ment_tco78 CLK_BASE->M2_ARSIZE[1]+3.161
pragma attribute SERDESIF_075 ment_tco79 CLK_BASE->M2_ARVALID+3.171
pragma attribute SERDESIF_075 ment_tco80 CLK_BASE->M2_AWADDR_HADDR[10]+3.057
pragma attribute SERDESIF_075 ment_tco81 CLK_BASE->M2_AWADDR_HADDR[11]+3.038
pragma attribute SERDESIF_075 ment_tco82 CLK_BASE->M2_AWADDR_HADDR[12]+3.093
pragma attribute SERDESIF_075 ment_tco83 CLK_BASE->M2_AWADDR_HADDR[13]+3.040
pragma attribute SERDESIF_075 ment_tco84 CLK_BASE->M2_AWADDR_HADDR[14]+3.051
pragma attribute SERDESIF_075 ment_tco85 CLK_BASE->M2_AWADDR_HADDR[15]+3.105
pragma attribute SERDESIF_075 ment_tco86 CLK_BASE->M2_AWADDR_HADDR[16]+3.087
pragma attribute SERDESIF_075 ment_tco87 CLK_BASE->M2_AWADDR_HADDR[17]+3.095
pragma attribute SERDESIF_075 ment_tco88 CLK_BASE->M2_AWADDR_HADDR[18]+3.123
pragma attribute SERDESIF_075 ment_tco89 CLK_BASE->M2_AWADDR_HADDR[19]+3.057
pragma attribute SERDESIF_075 ment_tco90 CLK_BASE->M2_AWADDR_HADDR[20]+3.167
pragma attribute SERDESIF_075 ment_tco91 CLK_BASE->M2_AWADDR_HADDR[21]+3.124
pragma attribute SERDESIF_075 ment_tco92 CLK_BASE->M2_AWADDR_HADDR[22]+3.054
pragma attribute SERDESIF_075 ment_tco93 CLK_BASE->M2_AWADDR_HADDR[23]+3.033
pragma attribute SERDESIF_075 ment_tco94 CLK_BASE->M2_AWADDR_HADDR[24]+3.125
pragma attribute SERDESIF_075 ment_tco95 CLK_BASE->M2_AWADDR_HADDR[25]+3.047
pragma attribute SERDESIF_075 ment_tco96 CLK_BASE->M2_AWADDR_HADDR[26]+3.076
pragma attribute SERDESIF_075 ment_tco97 CLK_BASE->M2_AWADDR_HADDR[27]+3.046
pragma attribute SERDESIF_075 ment_tco98 CLK_BASE->M2_AWADDR_HADDR[28]+3.058
pragma attribute SERDESIF_075 ment_tco99 CLK_BASE->M2_AWADDR_HADDR[29]+3.215
pragma attribute SERDESIF_075 ment_tco100 CLK_BASE->M2_AWADDR_HADDR[2]+3.132
pragma attribute SERDESIF_075 ment_tco101 CLK_BASE->M2_AWADDR_HADDR[30]+3.168
pragma attribute SERDESIF_075 ment_tco102 CLK_BASE->M2_AWADDR_HADDR[31]+3.035
pragma attribute SERDESIF_075 ment_tco103 CLK_BASE->M2_AWADDR_HADDR[3]+3.181
pragma attribute SERDESIF_075 ment_tco104 CLK_BASE->M2_AWADDR_HADDR[4]+3.044
pragma attribute SERDESIF_075 ment_tco105 CLK_BASE->M2_AWADDR_HADDR[5]+3.242
pragma attribute SERDESIF_075 ment_tco106 CLK_BASE->M2_AWADDR_HADDR[6]+3.248
pragma attribute SERDESIF_075 ment_tco107 CLK_BASE->M2_AWADDR_HADDR[7]+3.182
pragma attribute SERDESIF_075 ment_tco108 CLK_BASE->M2_AWADDR_HADDR[8]+3.239
pragma attribute SERDESIF_075 ment_tco109 CLK_BASE->M2_AWADDR_HADDR[9]+3.035
pragma attribute SERDESIF_075 ment_tco110 CLK_BASE->M2_AWBURST_HTRANS[0]+3.188
pragma attribute SERDESIF_075 ment_tco111 CLK_BASE->M2_AWLEN_HBURST[0]+3.007
pragma attribute SERDESIF_075 ment_tco112 CLK_BASE->M2_AWLEN_HBURST[1]+3.010
pragma attribute SERDESIF_075 ment_tco113 CLK_BASE->M2_AWLEN_HBURST[2]+3.006
pragma attribute SERDESIF_075 ment_tco114 CLK_BASE->M2_AWLEN_HBURST[3]+3.035
pragma attribute SERDESIF_075 ment_tco115 CLK_BASE->M2_AWSIZE_HSIZE[0]+3.064
pragma attribute SERDESIF_075 ment_tco116 CLK_BASE->M2_AWSIZE_HSIZE[1]+3.026
pragma attribute SERDESIF_075 ment_tco117 CLK_BASE->M2_AWVALID_HWRITE+3.190
pragma attribute SERDESIF_075 ment_tco118 CLK_BASE->M2_BREADY+3.185
pragma attribute SERDESIF_075 ment_tco119 CLK_BASE->M2_RREADY+2.845
pragma attribute SERDESIF_075 ment_tco120 CLK_BASE->M2_WDATA_HWDATA[0]+3.172
pragma attribute SERDESIF_075 ment_tco121 CLK_BASE->M2_WDATA_HWDATA[10]+3.234
pragma attribute SERDESIF_075 ment_tco122 CLK_BASE->M2_WDATA_HWDATA[11]+3.271
pragma attribute SERDESIF_075 ment_tco123 CLK_BASE->M2_WDATA_HWDATA[12]+3.269
pragma attribute SERDESIF_075 ment_tco124 CLK_BASE->M2_WDATA_HWDATA[13]+3.185
pragma attribute SERDESIF_075 ment_tco125 CLK_BASE->M2_WDATA_HWDATA[14]+3.244
pragma attribute SERDESIF_075 ment_tco126 CLK_BASE->M2_WDATA_HWDATA[15]+3.234
pragma attribute SERDESIF_075 ment_tco127 CLK_BASE->M2_WDATA_HWDATA[16]+3.248
pragma attribute SERDESIF_075 ment_tco128 CLK_BASE->M2_WDATA_HWDATA[17]+3.137
pragma attribute SERDESIF_075 ment_tco129 CLK_BASE->M2_WDATA_HWDATA[18]+3.193
pragma attribute SERDESIF_075 ment_tco130 CLK_BASE->M2_WDATA_HWDATA[19]+3.145
pragma attribute SERDESIF_075 ment_tco131 CLK_BASE->M2_WDATA_HWDATA[1]+3.150
pragma attribute SERDESIF_075 ment_tco132 CLK_BASE->M2_WDATA_HWDATA[20]+3.141
pragma attribute SERDESIF_075 ment_tco133 CLK_BASE->M2_WDATA_HWDATA[21]+3.190
pragma attribute SERDESIF_075 ment_tco134 CLK_BASE->M2_WDATA_HWDATA[22]+3.111
pragma attribute SERDESIF_075 ment_tco135 CLK_BASE->M2_WDATA_HWDATA[23]+3.109
pragma attribute SERDESIF_075 ment_tco136 CLK_BASE->M2_WDATA_HWDATA[24]+3.156
pragma attribute SERDESIF_075 ment_tco137 CLK_BASE->M2_WDATA_HWDATA[25]+3.176
pragma attribute SERDESIF_075 ment_tco138 CLK_BASE->M2_WDATA_HWDATA[26]+3.153
pragma attribute SERDESIF_075 ment_tco139 CLK_BASE->M2_WDATA_HWDATA[27]+3.146
pragma attribute SERDESIF_075 ment_tco140 CLK_BASE->M2_WDATA_HWDATA[28]+3.146
pragma attribute SERDESIF_075 ment_tco141 CLK_BASE->M2_WDATA_HWDATA[29]+3.250
pragma attribute SERDESIF_075 ment_tco142 CLK_BASE->M2_WDATA_HWDATA[2]+3.152
pragma attribute SERDESIF_075 ment_tco143 CLK_BASE->M2_WDATA_HWDATA[30]+3.199
pragma attribute SERDESIF_075 ment_tco144 CLK_BASE->M2_WDATA_HWDATA[31]+3.120
pragma attribute SERDESIF_075 ment_tco145 CLK_BASE->M2_WDATA_HWDATA[32]+3.163
pragma attribute SERDESIF_075 ment_tco146 CLK_BASE->M2_WDATA_HWDATA[33]+3.155
pragma attribute SERDESIF_075 ment_tco147 CLK_BASE->M2_WDATA_HWDATA[34]+3.148
pragma attribute SERDESIF_075 ment_tco148 CLK_BASE->M2_WDATA_HWDATA[35]+3.191
pragma attribute SERDESIF_075 ment_tco149 CLK_BASE->M2_WDATA_HWDATA[36]+3.093
pragma attribute SERDESIF_075 ment_tco150 CLK_BASE->M2_WDATA_HWDATA[37]+3.198
pragma attribute SERDESIF_075 ment_tco151 CLK_BASE->M2_WDATA_HWDATA[38]+3.195
pragma attribute SERDESIF_075 ment_tco152 CLK_BASE->M2_WDATA_HWDATA[39]+3.183
pragma attribute SERDESIF_075 ment_tco153 CLK_BASE->M2_WDATA_HWDATA[3]+3.197
pragma attribute SERDESIF_075 ment_tco154 CLK_BASE->M2_WDATA_HWDATA[40]+3.230
pragma attribute SERDESIF_075 ment_tco155 CLK_BASE->M2_WDATA_HWDATA[41]+3.093
pragma attribute SERDESIF_075 ment_tco156 CLK_BASE->M2_WDATA_HWDATA[42]+3.165
pragma attribute SERDESIF_075 ment_tco157 CLK_BASE->M2_WDATA_HWDATA[43]+3.219
pragma attribute SERDESIF_075 ment_tco158 CLK_BASE->M2_WDATA_HWDATA[44]+3.148
pragma attribute SERDESIF_075 ment_tco159 CLK_BASE->M2_WDATA_HWDATA[45]+3.183
pragma attribute SERDESIF_075 ment_tco160 CLK_BASE->M2_WDATA_HWDATA[46]+3.234
pragma attribute SERDESIF_075 ment_tco161 CLK_BASE->M2_WDATA_HWDATA[47]+3.108
pragma attribute SERDESIF_075 ment_tco162 CLK_BASE->M2_WDATA_HWDATA[48]+3.255
pragma attribute SERDESIF_075 ment_tco163 CLK_BASE->M2_WDATA_HWDATA[49]+3.150
pragma attribute SERDESIF_075 ment_tco164 CLK_BASE->M2_WDATA_HWDATA[4]+3.168
pragma attribute SERDESIF_075 ment_tco165 CLK_BASE->M2_WDATA_HWDATA[50]+3.163
pragma attribute SERDESIF_075 ment_tco166 CLK_BASE->M2_WDATA_HWDATA[51]+3.097
pragma attribute SERDESIF_075 ment_tco167 CLK_BASE->M2_WDATA_HWDATA[52]+3.070
pragma attribute SERDESIF_075 ment_tco168 CLK_BASE->M2_WDATA_HWDATA[53]+3.190
pragma attribute SERDESIF_075 ment_tco169 CLK_BASE->M2_WDATA_HWDATA[54]+3.206
pragma attribute SERDESIF_075 ment_tco170 CLK_BASE->M2_WDATA_HWDATA[55]+3.117
pragma attribute SERDESIF_075 ment_tco171 CLK_BASE->M2_WDATA_HWDATA[56]+3.193
pragma attribute SERDESIF_075 ment_tco172 CLK_BASE->M2_WDATA_HWDATA[57]+3.102
pragma attribute SERDESIF_075 ment_tco173 CLK_BASE->M2_WDATA_HWDATA[58]+3.073
pragma attribute SERDESIF_075 ment_tco174 CLK_BASE->M2_WDATA_HWDATA[59]+3.082
pragma attribute SERDESIF_075 ment_tco175 CLK_BASE->M2_WDATA_HWDATA[5]+3.139
pragma attribute SERDESIF_075 ment_tco176 CLK_BASE->M2_WDATA_HWDATA[60]+3.185
pragma attribute SERDESIF_075 ment_tco177 CLK_BASE->M2_WDATA_HWDATA[61]+3.144
pragma attribute SERDESIF_075 ment_tco178 CLK_BASE->M2_WDATA_HWDATA[62]+3.190
pragma attribute SERDESIF_075 ment_tco179 CLK_BASE->M2_WDATA_HWDATA[63]+3.145
pragma attribute SERDESIF_075 ment_tco180 CLK_BASE->M2_WDATA_HWDATA[6]+3.214
pragma attribute SERDESIF_075 ment_tco181 CLK_BASE->M2_WDATA_HWDATA[7]+3.172
pragma attribute SERDESIF_075 ment_tco182 CLK_BASE->M2_WDATA_HWDATA[8]+3.170
pragma attribute SERDESIF_075 ment_tco183 CLK_BASE->M2_WDATA_HWDATA[9]+3.104
pragma attribute SERDESIF_075 ment_tco184 CLK_BASE->M2_WLAST+3.097
pragma attribute SERDESIF_075 ment_tco185 CLK_BASE->M2_WSTRB[0]+3.174
pragma attribute SERDESIF_075 ment_tco186 CLK_BASE->M2_WSTRB[1]+3.168
pragma attribute SERDESIF_075 ment_tco187 CLK_BASE->M2_WSTRB[2]+3.249
pragma attribute SERDESIF_075 ment_tco188 CLK_BASE->M2_WSTRB[3]+3.145
pragma attribute SERDESIF_075 ment_tco189 CLK_BASE->M2_WSTRB[4]+3.294
pragma attribute SERDESIF_075 ment_tco190 CLK_BASE->M2_WSTRB[5]+3.129
pragma attribute SERDESIF_075 ment_tco191 CLK_BASE->M2_WSTRB[6]+3.172
pragma attribute SERDESIF_075 ment_tco192 CLK_BASE->M2_WSTRB[7]+3.080
pragma attribute SERDESIF_075 ment_tco193 CLK_BASE->M2_WVALID+3.207
pragma attribute SERDESIF_075 ment_tco194 CLK_BASE->M_ARADDR[0]+3.191
pragma attribute SERDESIF_075 ment_tco195 CLK_BASE->M_ARADDR[10]+3.072
pragma attribute SERDESIF_075 ment_tco196 CLK_BASE->M_ARADDR[11]+3.066
pragma attribute SERDESIF_075 ment_tco197 CLK_BASE->M_ARADDR[12]+3.025
pragma attribute SERDESIF_075 ment_tco198 CLK_BASE->M_ARADDR[13]+3.099
pragma attribute SERDESIF_075 ment_tco199 CLK_BASE->M_ARADDR[14]+3.006
pragma attribute SERDESIF_075 ment_tco200 CLK_BASE->M_ARADDR[15]+3.037
pragma attribute SERDESIF_075 ment_tco201 CLK_BASE->M_ARADDR[16]+3.112
pragma attribute SERDESIF_075 ment_tco202 CLK_BASE->M_ARADDR[17]+3.007
pragma attribute SERDESIF_075 ment_tco203 CLK_BASE->M_ARADDR[18]+3.168
pragma attribute SERDESIF_075 ment_tco204 CLK_BASE->M_ARADDR[19]+3.079
pragma attribute SERDESIF_075 ment_tco205 CLK_BASE->M_ARADDR[1]+3.211
pragma attribute SERDESIF_075 ment_tco206 CLK_BASE->M_ARADDR[20]+3.197
pragma attribute SERDESIF_075 ment_tco207 CLK_BASE->M_ARADDR[21]+3.144
pragma attribute SERDESIF_075 ment_tco208 CLK_BASE->M_ARADDR[22]+3.163
pragma attribute SERDESIF_075 ment_tco209 CLK_BASE->M_ARADDR[23]+3.196
pragma attribute SERDESIF_075 ment_tco210 CLK_BASE->M_ARADDR[24]+3.074
pragma attribute SERDESIF_075 ment_tco211 CLK_BASE->M_ARADDR[25]+3.147
pragma attribute SERDESIF_075 ment_tco212 CLK_BASE->M_ARADDR[26]+3.006
pragma attribute SERDESIF_075 ment_tco213 CLK_BASE->M_ARADDR[27]+2.989
pragma attribute SERDESIF_075 ment_tco214 CLK_BASE->M_ARADDR[28]+3.130
pragma attribute SERDESIF_075 ment_tco215 CLK_BASE->M_ARADDR[29]+3.033
pragma attribute SERDESIF_075 ment_tco216 CLK_BASE->M_ARADDR[2]+3.204
pragma attribute SERDESIF_075 ment_tco217 CLK_BASE->M_ARADDR[30]+3.071
pragma attribute SERDESIF_075 ment_tco218 CLK_BASE->M_ARADDR[31]+3.175
pragma attribute SERDESIF_075 ment_tco219 CLK_BASE->M_ARADDR[3]+3.195
pragma attribute SERDESIF_075 ment_tco220 CLK_BASE->M_ARADDR[4]+3.021
pragma attribute SERDESIF_075 ment_tco221 CLK_BASE->M_ARADDR[5]+3.038
pragma attribute SERDESIF_075 ment_tco222 CLK_BASE->M_ARADDR[6]+3.003
pragma attribute SERDESIF_075 ment_tco223 CLK_BASE->M_ARADDR[7]+3.061
pragma attribute SERDESIF_075 ment_tco224 CLK_BASE->M_ARADDR[8]+2.969
pragma attribute SERDESIF_075 ment_tco225 CLK_BASE->M_ARADDR[9]+3.015
pragma attribute SERDESIF_075 ment_tco226 CLK_BASE->M_ARBURST[0]+2.990
pragma attribute SERDESIF_075 ment_tco227 CLK_BASE->M_ARID[0]+2.933
pragma attribute SERDESIF_075 ment_tco228 CLK_BASE->M_ARID[1]+3.165
pragma attribute SERDESIF_075 ment_tco229 CLK_BASE->M_ARLEN[0]+2.909
pragma attribute SERDESIF_075 ment_tco230 CLK_BASE->M_ARLEN[1]+3.087
pragma attribute SERDESIF_075 ment_tco231 CLK_BASE->M_ARLEN[2]+3.050
pragma attribute SERDESIF_075 ment_tco232 CLK_BASE->M_ARLEN[3]+2.966
pragma attribute SERDESIF_075 ment_tco233 CLK_BASE->M_ARSIZE[0]+3.154
pragma attribute SERDESIF_075 ment_tco234 CLK_BASE->M_ARSIZE[1]+3.170
pragma attribute SERDESIF_075 ment_tco235 CLK_BASE->M_ARVALID+3.163
pragma attribute SERDESIF_075 ment_tco236 CLK_BASE->M_AWADDR_HADDR[10]+3.118
pragma attribute SERDESIF_075 ment_tco237 CLK_BASE->M_AWADDR_HADDR[11]+3.061
pragma attribute SERDESIF_075 ment_tco238 CLK_BASE->M_AWADDR_HADDR[12]+2.992
pragma attribute SERDESIF_075 ment_tco239 CLK_BASE->M_AWADDR_HADDR[13]+3.002
pragma attribute SERDESIF_075 ment_tco240 CLK_BASE->M_AWADDR_HADDR[14]+3.046
pragma attribute SERDESIF_075 ment_tco241 CLK_BASE->M_AWADDR_HADDR[15]+2.916
pragma attribute SERDESIF_075 ment_tco242 CLK_BASE->M_AWADDR_HADDR[16]+3.030
pragma attribute SERDESIF_075 ment_tco243 CLK_BASE->M_AWADDR_HADDR[17]+2.982
pragma attribute SERDESIF_075 ment_tco244 CLK_BASE->M_AWADDR_HADDR[18]+3.009
pragma attribute SERDESIF_075 ment_tco245 CLK_BASE->M_AWADDR_HADDR[19]+3.051
pragma attribute SERDESIF_075 ment_tco246 CLK_BASE->M_AWADDR_HADDR[20]+3.011
pragma attribute SERDESIF_075 ment_tco247 CLK_BASE->M_AWADDR_HADDR[21]+3.062
pragma attribute SERDESIF_075 ment_tco248 CLK_BASE->M_AWADDR_HADDR[22]+2.973
pragma attribute SERDESIF_075 ment_tco249 CLK_BASE->M_AWADDR_HADDR[23]+3.059
pragma attribute SERDESIF_075 ment_tco250 CLK_BASE->M_AWADDR_HADDR[24]+3.049
pragma attribute SERDESIF_075 ment_tco251 CLK_BASE->M_AWADDR_HADDR[25]+2.884
pragma attribute SERDESIF_075 ment_tco252 CLK_BASE->M_AWADDR_HADDR[26]+2.839
pragma attribute SERDESIF_075 ment_tco253 CLK_BASE->M_AWADDR_HADDR[27]+3.070
pragma attribute SERDESIF_075 ment_tco254 CLK_BASE->M_AWADDR_HADDR[28]+2.827
pragma attribute SERDESIF_075 ment_tco255 CLK_BASE->M_AWADDR_HADDR[29]+3.016
pragma attribute SERDESIF_075 ment_tco256 CLK_BASE->M_AWADDR_HADDR[2]+3.090
pragma attribute SERDESIF_075 ment_tco257 CLK_BASE->M_AWADDR_HADDR[30]+2.824
pragma attribute SERDESIF_075 ment_tco258 CLK_BASE->M_AWADDR_HADDR[31]+3.068
pragma attribute SERDESIF_075 ment_tco259 CLK_BASE->M_AWADDR_HADDR[3]+3.139
pragma attribute SERDESIF_075 ment_tco260 CLK_BASE->M_AWADDR_HADDR[4]+2.902
pragma attribute SERDESIF_075 ment_tco261 CLK_BASE->M_AWADDR_HADDR[5]+2.863
pragma attribute SERDESIF_075 ment_tco262 CLK_BASE->M_AWADDR_HADDR[6]+3.000
pragma attribute SERDESIF_075 ment_tco263 CLK_BASE->M_AWADDR_HADDR[7]+3.103
pragma attribute SERDESIF_075 ment_tco264 CLK_BASE->M_AWADDR_HADDR[8]+2.932
pragma attribute SERDESIF_075 ment_tco265 CLK_BASE->M_AWADDR_HADDR[9]+3.033
pragma attribute SERDESIF_075 ment_tco266 CLK_BASE->M_AWBURST_HTRANS[0]+2.946
pragma attribute SERDESIF_075 ment_tco267 CLK_BASE->M_AWLEN_HBURST[0]+3.046
pragma attribute SERDESIF_075 ment_tco268 CLK_BASE->M_AWLEN_HBURST[1]+3.008
pragma attribute SERDESIF_075 ment_tco269 CLK_BASE->M_AWLEN_HBURST[2]+2.848
pragma attribute SERDESIF_075 ment_tco270 CLK_BASE->M_AWLEN_HBURST[3]+2.964
pragma attribute SERDESIF_075 ment_tco271 CLK_BASE->M_AWSIZE_HSIZE[0]+3.026
pragma attribute SERDESIF_075 ment_tco272 CLK_BASE->M_AWSIZE_HSIZE[1]+2.902
pragma attribute SERDESIF_075 ment_tco273 CLK_BASE->M_AWVALID_HWRITE+3.046
pragma attribute SERDESIF_075 ment_tco274 CLK_BASE->M_BREADY+2.742
pragma attribute SERDESIF_075 ment_tco275 CLK_BASE->M_RREADY+3.100
pragma attribute SERDESIF_075 ment_tco276 CLK_BASE->M_WDATA_HWDATA[0]+3.746
pragma attribute SERDESIF_075 ment_tco277 CLK_BASE->M_WDATA_HWDATA[10]+4.000
pragma attribute SERDESIF_075 ment_tco278 CLK_BASE->M_WDATA_HWDATA[11]+3.531
pragma attribute SERDESIF_075 ment_tco279 CLK_BASE->M_WDATA_HWDATA[12]+3.870
pragma attribute SERDESIF_075 ment_tco280 CLK_BASE->M_WDATA_HWDATA[13]+3.741
pragma attribute SERDESIF_075 ment_tco281 CLK_BASE->M_WDATA_HWDATA[14]+3.770
pragma attribute SERDESIF_075 ment_tco282 CLK_BASE->M_WDATA_HWDATA[15]+3.868
pragma attribute SERDESIF_075 ment_tco283 CLK_BASE->M_WDATA_HWDATA[16]+3.822
pragma attribute SERDESIF_075 ment_tco284 CLK_BASE->M_WDATA_HWDATA[17]+3.808
pragma attribute SERDESIF_075 ment_tco285 CLK_BASE->M_WDATA_HWDATA[18]+3.574
pragma attribute SERDESIF_075 ment_tco286 CLK_BASE->M_WDATA_HWDATA[19]+3.982
pragma attribute SERDESIF_075 ment_tco287 CLK_BASE->M_WDATA_HWDATA[1]+3.500
pragma attribute SERDESIF_075 ment_tco288 CLK_BASE->M_WDATA_HWDATA[20]+3.893
pragma attribute SERDESIF_075 ment_tco289 CLK_BASE->M_WDATA_HWDATA[21]+3.755
pragma attribute SERDESIF_075 ment_tco290 CLK_BASE->M_WDATA_HWDATA[22]+3.780
pragma attribute SERDESIF_075 ment_tco291 CLK_BASE->M_WDATA_HWDATA[23]+3.517
pragma attribute SERDESIF_075 ment_tco292 CLK_BASE->M_WDATA_HWDATA[24]+3.710
pragma attribute SERDESIF_075 ment_tco293 CLK_BASE->M_WDATA_HWDATA[25]+3.607
pragma attribute SERDESIF_075 ment_tco294 CLK_BASE->M_WDATA_HWDATA[26]+3.583
pragma attribute SERDESIF_075 ment_tco295 CLK_BASE->M_WDATA_HWDATA[27]+3.540
pragma attribute SERDESIF_075 ment_tco296 CLK_BASE->M_WDATA_HWDATA[28]+3.547
pragma attribute SERDESIF_075 ment_tco297 CLK_BASE->M_WDATA_HWDATA[29]+3.697
pragma attribute SERDESIF_075 ment_tco298 CLK_BASE->M_WDATA_HWDATA[2]+3.859
pragma attribute SERDESIF_075 ment_tco299 CLK_BASE->M_WDATA_HWDATA[30]+3.528
pragma attribute SERDESIF_075 ment_tco300 CLK_BASE->M_WDATA_HWDATA[31]+3.316
pragma attribute SERDESIF_075 ment_tco301 CLK_BASE->M_WDATA_HWDATA[32]+3.433
pragma attribute SERDESIF_075 ment_tco302 CLK_BASE->M_WDATA_HWDATA[33]+3.408
pragma attribute SERDESIF_075 ment_tco303 CLK_BASE->M_WDATA_HWDATA[34]+3.210
pragma attribute SERDESIF_075 ment_tco304 CLK_BASE->M_WDATA_HWDATA[35]+3.448
pragma attribute SERDESIF_075 ment_tco305 CLK_BASE->M_WDATA_HWDATA[36]+3.297
pragma attribute SERDESIF_075 ment_tco306 CLK_BASE->M_WDATA_HWDATA[37]+3.214
pragma attribute SERDESIF_075 ment_tco307 CLK_BASE->M_WDATA_HWDATA[38]+3.290
pragma attribute SERDESIF_075 ment_tco308 CLK_BASE->M_WDATA_HWDATA[39]+3.256
pragma attribute SERDESIF_075 ment_tco309 CLK_BASE->M_WDATA_HWDATA[3]+3.869
pragma attribute SERDESIF_075 ment_tco310 CLK_BASE->M_WDATA_HWDATA[40]+3.252
pragma attribute SERDESIF_075 ment_tco311 CLK_BASE->M_WDATA_HWDATA[41]+3.362
pragma attribute SERDESIF_075 ment_tco312 CLK_BASE->M_WDATA_HWDATA[42]+3.435
pragma attribute SERDESIF_075 ment_tco313 CLK_BASE->M_WDATA_HWDATA[43]+3.448
pragma attribute SERDESIF_075 ment_tco314 CLK_BASE->M_WDATA_HWDATA[44]+3.283
pragma attribute SERDESIF_075 ment_tco315 CLK_BASE->M_WDATA_HWDATA[45]+3.458
pragma attribute SERDESIF_075 ment_tco316 CLK_BASE->M_WDATA_HWDATA[46]+3.312
pragma attribute SERDESIF_075 ment_tco317 CLK_BASE->M_WDATA_HWDATA[47]+3.530
pragma attribute SERDESIF_075 ment_tco318 CLK_BASE->M_WDATA_HWDATA[48]+3.379
pragma attribute SERDESIF_075 ment_tco319 CLK_BASE->M_WDATA_HWDATA[49]+3.323
pragma attribute SERDESIF_075 ment_tco320 CLK_BASE->M_WDATA_HWDATA[4]+3.846
pragma attribute SERDESIF_075 ment_tco321 CLK_BASE->M_WDATA_HWDATA[50]+3.320
pragma attribute SERDESIF_075 ment_tco322 CLK_BASE->M_WDATA_HWDATA[51]+3.452
pragma attribute SERDESIF_075 ment_tco323 CLK_BASE->M_WDATA_HWDATA[52]+3.666
pragma attribute SERDESIF_075 ment_tco324 CLK_BASE->M_WDATA_HWDATA[53]+3.846
pragma attribute SERDESIF_075 ment_tco325 CLK_BASE->M_WDATA_HWDATA[54]+3.682
pragma attribute SERDESIF_075 ment_tco326 CLK_BASE->M_WDATA_HWDATA[55]+3.489
pragma attribute SERDESIF_075 ment_tco327 CLK_BASE->M_WDATA_HWDATA[56]+3.628
pragma attribute SERDESIF_075 ment_tco328 CLK_BASE->M_WDATA_HWDATA[57]+3.583
pragma attribute SERDESIF_075 ment_tco329 CLK_BASE->M_WDATA_HWDATA[58]+3.502
pragma attribute SERDESIF_075 ment_tco330 CLK_BASE->M_WDATA_HWDATA[59]+3.729
pragma attribute SERDESIF_075 ment_tco331 CLK_BASE->M_WDATA_HWDATA[5]+3.708
pragma attribute SERDESIF_075 ment_tco332 CLK_BASE->M_WDATA_HWDATA[60]+3.535
pragma attribute SERDESIF_075 ment_tco333 CLK_BASE->M_WDATA_HWDATA[61]+3.626
pragma attribute SERDESIF_075 ment_tco334 CLK_BASE->M_WDATA_HWDATA[62]+3.781
pragma attribute SERDESIF_075 ment_tco335 CLK_BASE->M_WDATA_HWDATA[63]+3.621
pragma attribute SERDESIF_075 ment_tco336 CLK_BASE->M_WDATA_HWDATA[6]+3.684
pragma attribute SERDESIF_075 ment_tco337 CLK_BASE->M_WDATA_HWDATA[7]+3.796
pragma attribute SERDESIF_075 ment_tco338 CLK_BASE->M_WDATA_HWDATA[8]+3.568
pragma attribute SERDESIF_075 ment_tco339 CLK_BASE->M_WDATA_HWDATA[9]+3.651
pragma attribute SERDESIF_075 ment_tco340 CLK_BASE->M_WLAST+3.108
pragma attribute SERDESIF_075 ment_tco341 CLK_BASE->M_WSTRB[0]+3.237
pragma attribute SERDESIF_075 ment_tco342 CLK_BASE->M_WSTRB[1]+3.676
pragma attribute SERDESIF_075 ment_tco343 CLK_BASE->M_WSTRB[2]+3.572
pragma attribute SERDESIF_075 ment_tco344 CLK_BASE->M_WSTRB[3]+3.481
pragma attribute SERDESIF_075 ment_tco345 CLK_BASE->M_WSTRB[4]+3.574
pragma attribute SERDESIF_075 ment_tco346 CLK_BASE->M_WSTRB[5]+3.608
pragma attribute SERDESIF_075 ment_tco347 CLK_BASE->M_WSTRB[6]+3.429
pragma attribute SERDESIF_075 ment_tco348 CLK_BASE->M_WSTRB[7]+3.575
pragma attribute SERDESIF_075 ment_tco349 CLK_BASE->M_WVALID+3.090
pragma attribute SERDESIF_075 ment_tco350 CLK_BASE->S2_ARREADY+3.099
pragma attribute SERDESIF_075 ment_tco351 CLK_BASE->S2_AWREADY+3.067
pragma attribute SERDESIF_075 ment_tco352 CLK_BASE->S2_BID[0]+3.109
pragma attribute SERDESIF_075 ment_tco353 CLK_BASE->S2_BID[1]+3.104
pragma attribute SERDESIF_075 ment_tco354 CLK_BASE->S2_BID[2]+3.086
pragma attribute SERDESIF_075 ment_tco355 CLK_BASE->S2_BID[3]+3.045
pragma attribute SERDESIF_075 ment_tco356 CLK_BASE->S2_BRESP_HRESP[1]+3.194
pragma attribute SERDESIF_075 ment_tco357 CLK_BASE->S2_BVALID+3.152
pragma attribute SERDESIF_075 ment_tco358 CLK_BASE->S2_RDATA_HRDATA[0]+3.001
pragma attribute SERDESIF_075 ment_tco359 CLK_BASE->S2_RDATA_HRDATA[10]+3.047
pragma attribute SERDESIF_075 ment_tco360 CLK_BASE->S2_RDATA_HRDATA[11]+3.066
pragma attribute SERDESIF_075 ment_tco361 CLK_BASE->S2_RDATA_HRDATA[12]+3.070
pragma attribute SERDESIF_075 ment_tco362 CLK_BASE->S2_RDATA_HRDATA[13]+3.017
pragma attribute SERDESIF_075 ment_tco363 CLK_BASE->S2_RDATA_HRDATA[14]+3.034
pragma attribute SERDESIF_075 ment_tco364 CLK_BASE->S2_RDATA_HRDATA[15]+3.016
pragma attribute SERDESIF_075 ment_tco365 CLK_BASE->S2_RDATA_HRDATA[16]+3.039
pragma attribute SERDESIF_075 ment_tco366 CLK_BASE->S2_RDATA_HRDATA[17]+3.015
pragma attribute SERDESIF_075 ment_tco367 CLK_BASE->S2_RDATA_HRDATA[18]+3.000
pragma attribute SERDESIF_075 ment_tco368 CLK_BASE->S2_RDATA_HRDATA[19]+3.023
pragma attribute SERDESIF_075 ment_tco369 CLK_BASE->S2_RDATA_HRDATA[1]+2.991
pragma attribute SERDESIF_075 ment_tco370 CLK_BASE->S2_RDATA_HRDATA[20]+3.045
pragma attribute SERDESIF_075 ment_tco371 CLK_BASE->S2_RDATA_HRDATA[21]+3.006
pragma attribute SERDESIF_075 ment_tco372 CLK_BASE->S2_RDATA_HRDATA[22]+3.019
pragma attribute SERDESIF_075 ment_tco373 CLK_BASE->S2_RDATA_HRDATA[23]+3.014
pragma attribute SERDESIF_075 ment_tco374 CLK_BASE->S2_RDATA_HRDATA[24]+3.018
pragma attribute SERDESIF_075 ment_tco375 CLK_BASE->S2_RDATA_HRDATA[25]+3.058
pragma attribute SERDESIF_075 ment_tco376 CLK_BASE->S2_RDATA_HRDATA[26]+3.003
pragma attribute SERDESIF_075 ment_tco377 CLK_BASE->S2_RDATA_HRDATA[27]+3.108
pragma attribute SERDESIF_075 ment_tco378 CLK_BASE->S2_RDATA_HRDATA[28]+3.010
pragma attribute SERDESIF_075 ment_tco379 CLK_BASE->S2_RDATA_HRDATA[29]+2.980
pragma attribute SERDESIF_075 ment_tco380 CLK_BASE->S2_RDATA_HRDATA[2]+2.986
pragma attribute SERDESIF_075 ment_tco381 CLK_BASE->S2_RDATA_HRDATA[30]+2.964
pragma attribute SERDESIF_075 ment_tco382 CLK_BASE->S2_RDATA_HRDATA[31]+3.098
pragma attribute SERDESIF_075 ment_tco383 CLK_BASE->S2_RDATA_HRDATA[32]+3.044
pragma attribute SERDESIF_075 ment_tco384 CLK_BASE->S2_RDATA_HRDATA[33]+3.175
pragma attribute SERDESIF_075 ment_tco385 CLK_BASE->S2_RDATA_HRDATA[34]+3.131
pragma attribute SERDESIF_075 ment_tco386 CLK_BASE->S2_RDATA_HRDATA[35]+3.105
pragma attribute SERDESIF_075 ment_tco387 CLK_BASE->S2_RDATA_HRDATA[36]+3.146
pragma attribute SERDESIF_075 ment_tco388 CLK_BASE->S2_RDATA_HRDATA[37]+3.101
pragma attribute SERDESIF_075 ment_tco389 CLK_BASE->S2_RDATA_HRDATA[38]+3.026
pragma attribute SERDESIF_075 ment_tco390 CLK_BASE->S2_RDATA_HRDATA[39]+3.134
pragma attribute SERDESIF_075 ment_tco391 CLK_BASE->S2_RDATA_HRDATA[3]+2.967
pragma attribute SERDESIF_075 ment_tco392 CLK_BASE->S2_RDATA_HRDATA[40]+3.147
pragma attribute SERDESIF_075 ment_tco393 CLK_BASE->S2_RDATA_HRDATA[41]+3.089
pragma attribute SERDESIF_075 ment_tco394 CLK_BASE->S2_RDATA_HRDATA[42]+3.145
pragma attribute SERDESIF_075 ment_tco395 CLK_BASE->S2_RDATA_HRDATA[43]+3.139
pragma attribute SERDESIF_075 ment_tco396 CLK_BASE->S2_RDATA_HRDATA[44]+3.086
pragma attribute SERDESIF_075 ment_tco397 CLK_BASE->S2_RDATA_HRDATA[45]+3.174
pragma attribute SERDESIF_075 ment_tco398 CLK_BASE->S2_RDATA_HRDATA[46]+3.178
pragma attribute SERDESIF_075 ment_tco399 CLK_BASE->S2_RDATA_HRDATA[47]+3.119
pragma attribute SERDESIF_075 ment_tco400 CLK_BASE->S2_RDATA_HRDATA[48]+3.172
pragma attribute SERDESIF_075 ment_tco401 CLK_BASE->S2_RDATA_HRDATA[49]+3.060
pragma attribute SERDESIF_075 ment_tco402 CLK_BASE->S2_RDATA_HRDATA[4]+3.052
pragma attribute SERDESIF_075 ment_tco403 CLK_BASE->S2_RDATA_HRDATA[50]+3.157
pragma attribute SERDESIF_075 ment_tco404 CLK_BASE->S2_RDATA_HRDATA[51]+3.117
pragma attribute SERDESIF_075 ment_tco405 CLK_BASE->S2_RDATA_HRDATA[52]+3.175
pragma attribute SERDESIF_075 ment_tco406 CLK_BASE->S2_RDATA_HRDATA[53]+3.053
pragma attribute SERDESIF_075 ment_tco407 CLK_BASE->S2_RDATA_HRDATA[54]+3.111
pragma attribute SERDESIF_075 ment_tco408 CLK_BASE->S2_RDATA_HRDATA[55]+3.064
pragma attribute SERDESIF_075 ment_tco409 CLK_BASE->S2_RDATA_HRDATA[56]+3.159
pragma attribute SERDESIF_075 ment_tco410 CLK_BASE->S2_RDATA_HRDATA[57]+3.093
pragma attribute SERDESIF_075 ment_tco411 CLK_BASE->S2_RDATA_HRDATA[58]+3.150
pragma attribute SERDESIF_075 ment_tco412 CLK_BASE->S2_RDATA_HRDATA[59]+3.088
pragma attribute SERDESIF_075 ment_tco413 CLK_BASE->S2_RDATA_HRDATA[5]+3.082
pragma attribute SERDESIF_075 ment_tco414 CLK_BASE->S2_RDATA_HRDATA[60]+3.101
pragma attribute SERDESIF_075 ment_tco415 CLK_BASE->S2_RDATA_HRDATA[61]+3.029
pragma attribute SERDESIF_075 ment_tco416 CLK_BASE->S2_RDATA_HRDATA[62]+2.968
pragma attribute SERDESIF_075 ment_tco417 CLK_BASE->S2_RDATA_HRDATA[63]+3.044
pragma attribute SERDESIF_075 ment_tco418 CLK_BASE->S2_RDATA_HRDATA[6]+3.065
pragma attribute SERDESIF_075 ment_tco419 CLK_BASE->S2_RDATA_HRDATA[7]+3.012
pragma attribute SERDESIF_075 ment_tco420 CLK_BASE->S2_RDATA_HRDATA[8]+3.036
pragma attribute SERDESIF_075 ment_tco421 CLK_BASE->S2_RDATA_HRDATA[9]+3.005
pragma attribute SERDESIF_075 ment_tco422 CLK_BASE->S2_RID[0]+2.927
pragma attribute SERDESIF_075 ment_tco423 CLK_BASE->S2_RID[1]+3.011
pragma attribute SERDESIF_075 ment_tco424 CLK_BASE->S2_RID[2]+3.018
pragma attribute SERDESIF_075 ment_tco425 CLK_BASE->S2_RID[3]+2.942
pragma attribute SERDESIF_075 ment_tco426 CLK_BASE->S2_RLAST+3.084
pragma attribute SERDESIF_075 ment_tco427 CLK_BASE->S2_RRESP[1]+2.948
pragma attribute SERDESIF_075 ment_tco428 CLK_BASE->S2_RVALID+3.161
pragma attribute SERDESIF_075 ment_tco429 CLK_BASE->S2_WREADY_HREADYOUT+2.645
pragma attribute SERDESIF_075 ment_tco430 CLK_BASE->S_ARREADY+2.901
pragma attribute SERDESIF_075 ment_tco431 CLK_BASE->S_AWREADY+2.934
pragma attribute SERDESIF_075 ment_tco432 CLK_BASE->S_BID[0]+3.098
pragma attribute SERDESIF_075 ment_tco433 CLK_BASE->S_BID[1]+3.147
pragma attribute SERDESIF_075 ment_tco434 CLK_BASE->S_BID[2]+3.169
pragma attribute SERDESIF_075 ment_tco435 CLK_BASE->S_BID[3]+3.215
pragma attribute SERDESIF_075 ment_tco436 CLK_BASE->S_BRESP_HRESP[1]+3.199
pragma attribute SERDESIF_075 ment_tco437 CLK_BASE->S_BVALID+3.251
pragma attribute SERDESIF_075 ment_tco438 CLK_BASE->S_RDATA_HRDATA[0]+3.170
pragma attribute SERDESIF_075 ment_tco439 CLK_BASE->S_RDATA_HRDATA[10]+3.148
pragma attribute SERDESIF_075 ment_tco440 CLK_BASE->S_RDATA_HRDATA[11]+3.170
pragma attribute SERDESIF_075 ment_tco441 CLK_BASE->S_RDATA_HRDATA[12]+3.164
pragma attribute SERDESIF_075 ment_tco442 CLK_BASE->S_RDATA_HRDATA[13]+3.137
pragma attribute SERDESIF_075 ment_tco443 CLK_BASE->S_RDATA_HRDATA[14]+3.161
pragma attribute SERDESIF_075 ment_tco444 CLK_BASE->S_RDATA_HRDATA[15]+3.150
pragma attribute SERDESIF_075 ment_tco445 CLK_BASE->S_RDATA_HRDATA[16]+3.186
pragma attribute SERDESIF_075 ment_tco446 CLK_BASE->S_RDATA_HRDATA[17]+3.128
pragma attribute SERDESIF_075 ment_tco447 CLK_BASE->S_RDATA_HRDATA[18]+3.142
pragma attribute SERDESIF_075 ment_tco448 CLK_BASE->S_RDATA_HRDATA[19]+3.181
pragma attribute SERDESIF_075 ment_tco449 CLK_BASE->S_RDATA_HRDATA[1]+3.155
pragma attribute SERDESIF_075 ment_tco450 CLK_BASE->S_RDATA_HRDATA[20]+3.159
pragma attribute SERDESIF_075 ment_tco451 CLK_BASE->S_RDATA_HRDATA[21]+3.128
pragma attribute SERDESIF_075 ment_tco452 CLK_BASE->S_RDATA_HRDATA[22]+3.146
pragma attribute SERDESIF_075 ment_tco453 CLK_BASE->S_RDATA_HRDATA[23]+3.170
pragma attribute SERDESIF_075 ment_tco454 CLK_BASE->S_RDATA_HRDATA[24]+3.185
pragma attribute SERDESIF_075 ment_tco455 CLK_BASE->S_RDATA_HRDATA[25]+3.220
pragma attribute SERDESIF_075 ment_tco456 CLK_BASE->S_RDATA_HRDATA[26]+3.180
pragma attribute SERDESIF_075 ment_tco457 CLK_BASE->S_RDATA_HRDATA[27]+3.188
pragma attribute SERDESIF_075 ment_tco458 CLK_BASE->S_RDATA_HRDATA[28]+3.141
pragma attribute SERDESIF_075 ment_tco459 CLK_BASE->S_RDATA_HRDATA[29]+3.175
pragma attribute SERDESIF_075 ment_tco460 CLK_BASE->S_RDATA_HRDATA[2]+3.139
pragma attribute SERDESIF_075 ment_tco461 CLK_BASE->S_RDATA_HRDATA[30]+3.170
pragma attribute SERDESIF_075 ment_tco462 CLK_BASE->S_RDATA_HRDATA[31]+3.183
pragma attribute SERDESIF_075 ment_tco463 CLK_BASE->S_RDATA_HRDATA[32]+3.285
pragma attribute SERDESIF_075 ment_tco464 CLK_BASE->S_RDATA_HRDATA[33]+3.299
pragma attribute SERDESIF_075 ment_tco465 CLK_BASE->S_RDATA_HRDATA[34]+3.362
pragma attribute SERDESIF_075 ment_tco466 CLK_BASE->S_RDATA_HRDATA[35]+3.306
pragma attribute SERDESIF_075 ment_tco467 CLK_BASE->S_RDATA_HRDATA[36]+3.256
pragma attribute SERDESIF_075 ment_tco468 CLK_BASE->S_RDATA_HRDATA[37]+3.260
pragma attribute SERDESIF_075 ment_tco469 CLK_BASE->S_RDATA_HRDATA[38]+3.263
pragma attribute SERDESIF_075 ment_tco470 CLK_BASE->S_RDATA_HRDATA[39]+3.294
pragma attribute SERDESIF_075 ment_tco471 CLK_BASE->S_RDATA_HRDATA[3]+3.178
pragma attribute SERDESIF_075 ment_tco472 CLK_BASE->S_RDATA_HRDATA[40]+3.277
pragma attribute SERDESIF_075 ment_tco473 CLK_BASE->S_RDATA_HRDATA[41]+3.293
pragma attribute SERDESIF_075 ment_tco474 CLK_BASE->S_RDATA_HRDATA[42]+3.261
pragma attribute SERDESIF_075 ment_tco475 CLK_BASE->S_RDATA_HRDATA[43]+3.304
pragma attribute SERDESIF_075 ment_tco476 CLK_BASE->S_RDATA_HRDATA[44]+3.432
pragma attribute SERDESIF_075 ment_tco477 CLK_BASE->S_RDATA_HRDATA[45]+3.389
pragma attribute SERDESIF_075 ment_tco478 CLK_BASE->S_RDATA_HRDATA[46]+3.439
pragma attribute SERDESIF_075 ment_tco479 CLK_BASE->S_RDATA_HRDATA[47]+3.312
pragma attribute SERDESIF_075 ment_tco480 CLK_BASE->S_RDATA_HRDATA[48]+3.284
pragma attribute SERDESIF_075 ment_tco481 CLK_BASE->S_RDATA_HRDATA[49]+3.246
pragma attribute SERDESIF_075 ment_tco482 CLK_BASE->S_RDATA_HRDATA[4]+3.132
pragma attribute SERDESIF_075 ment_tco483 CLK_BASE->S_RDATA_HRDATA[50]+3.289
pragma attribute SERDESIF_075 ment_tco484 CLK_BASE->S_RDATA_HRDATA[51]+3.233
pragma attribute SERDESIF_075 ment_tco485 CLK_BASE->S_RDATA_HRDATA[52]+3.175
pragma attribute SERDESIF_075 ment_tco486 CLK_BASE->S_RDATA_HRDATA[53]+3.163
pragma attribute SERDESIF_075 ment_tco487 CLK_BASE->S_RDATA_HRDATA[54]+3.157
pragma attribute SERDESIF_075 ment_tco488 CLK_BASE->S_RDATA_HRDATA[55]+3.169
pragma attribute SERDESIF_075 ment_tco489 CLK_BASE->S_RDATA_HRDATA[56]+3.169
pragma attribute SERDESIF_075 ment_tco490 CLK_BASE->S_RDATA_HRDATA[57]+3.147
pragma attribute SERDESIF_075 ment_tco491 CLK_BASE->S_RDATA_HRDATA[58]+3.140
pragma attribute SERDESIF_075 ment_tco492 CLK_BASE->S_RDATA_HRDATA[59]+3.196
pragma attribute SERDESIF_075 ment_tco493 CLK_BASE->S_RDATA_HRDATA[5]+3.126
pragma attribute SERDESIF_075 ment_tco494 CLK_BASE->S_RDATA_HRDATA[60]+3.181
pragma attribute SERDESIF_075 ment_tco495 CLK_BASE->S_RDATA_HRDATA[61]+3.210
pragma attribute SERDESIF_075 ment_tco496 CLK_BASE->S_RDATA_HRDATA[62]+3.199
pragma attribute SERDESIF_075 ment_tco497 CLK_BASE->S_RDATA_HRDATA[63]+3.143
pragma attribute SERDESIF_075 ment_tco498 CLK_BASE->S_RDATA_HRDATA[6]+3.176
pragma attribute SERDESIF_075 ment_tco499 CLK_BASE->S_RDATA_HRDATA[7]+3.169
pragma attribute SERDESIF_075 ment_tco500 CLK_BASE->S_RDATA_HRDATA[8]+3.209
pragma attribute SERDESIF_075 ment_tco501 CLK_BASE->S_RDATA_HRDATA[9]+3.125
pragma attribute SERDESIF_075 ment_tco502 CLK_BASE->S_RID[0]+3.275
pragma attribute SERDESIF_075 ment_tco503 CLK_BASE->S_RID[1]+3.215
pragma attribute SERDESIF_075 ment_tco504 CLK_BASE->S_RID[2]+3.140
pragma attribute SERDESIF_075 ment_tco505 CLK_BASE->S_RID[3]+3.162
pragma attribute SERDESIF_075 ment_tco506 CLK_BASE->S_RLAST+3.242
pragma attribute SERDESIF_075 ment_tco507 CLK_BASE->S_RRESP[1]+3.150
pragma attribute SERDESIF_075 ment_tco508 CLK_BASE->S_RVALID+3.122
pragma attribute SERDESIF_075 ment_tco509 CLK_BASE->S_WREADY_HREADYOUT+2.805
*/
/* synthesis black_box black_box_pad ="RXD3_P,RXD2_P,RXD1_P,RXD0_P,RXD3_N,RXD2_N,RXD1_N,RXD0_N,TXD3_P,TXD2_P,TXD1_P,TXD0_P,TXD3_N,TXD2_N,TXD1_N,TXD0_N" */
 ;
output [31:0] APB_PRDATA;
output APB_PREADY;
output APB_PSLVERR;
output [1:0] ATXCLKSTABLE;
output [1:0] EPCS_READY;
output [1:0] EPCS_RXCLK;
output EPCS_RXCLK_0;
output EPCS_RXCLK_1;
output [39:0] EPCS_RXDATA;
output [1:0] EPCS_RXIDLE;
output [1:0] EPCS_RXRSTN;
output [1:0] EPCS_RXVAL;
output [1:0] EPCS_TXCLK;
output EPCS_TXCLK_0;
output EPCS_TXCLK_1;
output [1:0] EPCS_TXRSTN;
output FATC_RESET_N;
output H2FCALIB0;
output H2FCALIB1;
output [31:0] M2_ARADDR;
output [1:0] M2_ARBURST;
output [3:0] M2_ARID;
output [3:0] M2_ARLEN;
output [1:0] M2_ARSIZE;
output M2_ARVALID;
output [31:0] M2_AWADDR_HADDR;
output [1:0] M2_AWBURST_HTRANS;
output [3:0] M2_AWID;
output [3:0] M2_AWLEN_HBURST;
output [1:0] M2_AWSIZE_HSIZE;
output M2_AWVALID_HWRITE;
output M2_BREADY;
output M2_RREADY;
output [63:0] M2_WDATA_HWDATA;
output [3:0] M2_WID;
output M2_WLAST;
output [7:0] M2_WSTRB;
output M2_WVALID;
output [31:0] M_ARADDR;
output [1:0] M_ARBURST;
output [3:0] M_ARID;
output [3:0] M_ARLEN;
output [1:0] M_ARSIZE;
output M_ARVALID;
output [31:0] M_AWADDR_HADDR;
output [1:0] M_AWBURST_HTRANS;
output [3:0] M_AWID;
output [3:0] M_AWLEN_HBURST;
output [1:0] M_AWSIZE_HSIZE;
output M_AWVALID_HWRITE;
output M_BREADY;
output M_RREADY;
output [63:0] M_WDATA_HWDATA;
output [3:0] M_WID;
output M_WLAST;
output [7:0] M_WSTRB;
output M_WVALID;
output [5:0] PCIE2_LTSSM;
output PCIE2_SYSTEM_INT;
output PCIE2_WAKE_N;
output [5:0] PCIE_LTSSM;
output PCIE_SYSTEM_INT;
output PLL_LOCK_INT;
output PLL_LOCKLOST_INT;
output S2_ARREADY;
output S2_AWREADY;
output [3:0] S2_BID;
output [1:0] S2_BRESP_HRESP;
output S2_BVALID;
output [63:0] S2_RDATA_HRDATA;
output [3:0] S2_RID;
output S2_RLAST;
output [1:0] S2_RRESP;
output S2_RVALID;
output S2_WREADY_HREADYOUT;
output S_ARREADY;
output S_AWREADY;
output [3:0] S_BID;
output [1:0] S_BRESP_HRESP;
output S_BVALID;
output [63:0] S_RDATA_HRDATA;
output [3:0] S_RID;
output S_RLAST;
output [1:0] S_RRESP;
output S_RVALID;
output S_WREADY_HREADYOUT;
output SPLL_LOCK;
output WAKE_N;
output XAUI_OUT_CLK;
input  APB_CLK;
input  [14:2] APB_PADDR;
input  APB_PENABLE;
input  APB_PSEL;
input  [31:0] APB_PWDATA;
input  APB_PWRITE;
input  APB_RSTN;
input  CLK_BASE;
input  [1:0] EPCS_PWRDN;
input  [1:0] EPCS_RSTN;
input  [1:0] EPCS_RXERR;
input  [39:0] EPCS_TXDATA;
input  [1:0] EPCS_TXOOB;
input  [1:0] EPCS_TXVAL;
input  F2HCALIB0;
input  F2HCALIB1;
input  FAB_PLL_LOCK;
input  FAB_REF_CLK;
input  M2_ARREADY;
input  M2_AWREADY;
input  [3:0] M2_BID;
input  [1:0] M2_BRESP_HRESP;
input  M2_BVALID;
input  [63:0] M2_RDATA_HRDATA;
input  [3:0] M2_RID;
input  M2_RLAST;
input  [1:0] M2_RRESP;
input  M2_RVALID;
input  M2_WREADY_HREADY;
input  M_ARREADY;
input  M_AWREADY;
input  [3:0] M_BID;
input  [1:0] M_BRESP_HRESP;
input  M_BVALID;
input  [63:0] M_RDATA_HRDATA;
input  [3:0] M_RID;
input  M_RLAST;
input  [1:0] M_RRESP;
input  M_RVALID;
input  M_WREADY_HREADY;
input  [3:0] PCIE2_INTERRUPT;
input  PCIE2_PERST_N;
input  PCIE2_SERDESIF_CORE_RESET_N;
input  PCIE2_WAKE_REQ;
input  [3:0] PCIE_INTERRUPT;
input  PERST_N;
input  [31:0] S2_ARADDR;
input  [1:0] S2_ARBURST;
input  [3:0] S2_ARID;
input  [3:0] S2_ARLEN;
input  [1:0] S2_ARLOCK;
input  [1:0] S2_ARSIZE;
input  S2_ARVALID;
input  [31:0] S2_AWADDR_HADDR;
input  [1:0] S2_AWBURST_HTRANS;
input  [3:0] S2_AWID_HSEL;
input  [3:0] S2_AWLEN_HBURST;
input  [1:0] S2_AWLOCK;
input  [1:0] S2_AWSIZE_HSIZE;
input  S2_AWVALID_HWRITE;
input  S2_BREADY_HREADY;
input  S2_RREADY;
input  [63:0] S2_WDATA_HWDATA;
input  [3:0] S2_WID;
input  S2_WLAST;
input  [7:0] S2_WSTRB;
input  S2_WVALID;
input  [31:0] S_ARADDR;
input  [1:0] S_ARBURST;
input  [3:0] S_ARID;
input  [3:0] S_ARLEN;
input  [1:0] S_ARLOCK;
input  [1:0] S_ARSIZE;
input  S_ARVALID;
input  [31:0] S_AWADDR_HADDR;
input  [1:0] S_AWBURST_HTRANS;
input  [3:0] S_AWID_HSEL;
input  [3:0] S_AWLEN_HBURST;
input  [1:0] S_AWLOCK;
input  [1:0] S_AWSIZE_HSIZE;
input  S_AWVALID_HWRITE;
input  S_BREADY_HREADY;
input  S_RREADY;
input  [63:0] S_WDATA_HWDATA;
input  [3:0] S_WID;
input  S_WLAST;
input  [7:0] S_WSTRB;
input  S_WVALID;
input  SERDESIF_CORE_RESET_N;
input  SERDESIF_PHY_RESET_N;
input  WAKE_REQ;
input  XAUI_FB_CLK;
input  RXD3_P;
input  RXD2_P;
input  RXD1_P;
input  RXD0_P;
input  RXD3_N;
input  RXD2_N;
input  RXD1_N;
input  RXD0_N;
output TXD3_P;
output TXD2_P;
output TXD1_P;
output TXD0_P;
output TXD3_N;
output TXD2_N;
output TXD1_N;
output TXD0_N;
input  REFCLK0;
input  REFCLK1;
parameter INIT = 'h0;
parameter ACT_CONFIG = "";
parameter ACT_SIM = 0;

endmodule
